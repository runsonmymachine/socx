    bins HwsRomNetInit                                            = { [ (('h4000fc00 - 'h4000fc00) >> 1) : ((('h4000fc00 - 'h4000fc00 + 'd18) >> 1) - 1) ] };
    bins HwsRomFlowFSMPowerupB2B                                  = { [ (('h4000fc12 - 'h4000fc00) >> 1) : ((('h4000fc12 - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomFlowManagerOverlayInitFromGnvm                     = { [ (('h4000fc1a - 'h4000fc00) >> 1) : ((('h4000fc1a - 'h4000fc00 + 'd6) >> 1) - 1) ] };
    bins HwsRomTempSensingOverlayInitFromGnvm                     = { [ (('h4000fc20 - 'h4000fc00) >> 1) : ((('h4000fc20 - 'h4000fc00 + 'd6) >> 1) - 1) ] };
    bins HwsRomRxSweepAndAuxMeasOverlayInitFromGnvm               = { [ (('h4000fc26 - 'h4000fc00) >> 1) : ((('h4000fc26 - 'h4000fc00 + 'd6) >> 1) - 1) ] };
    bins HwsRomTempSenseLvRadioInit                               = { [ (('h4000fc2c - 'h4000fc00) >> 1) : ((('h4000fc2c - 'h4000fc00 + 'd14) >> 1) - 1) ] };
    bins HwsRomTempSenseLvActivation                              = { [ (('h4000fc3a - 'h4000fc00) >> 1) : ((('h4000fc3a - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomTempSensePopulateOvlB2B                            = { [ (('h4000fc42 - 'h4000fc00) >> 1) : ((('h4000fc42 - 'h4000fc00 + 'd4) >> 1) - 1) ] };
    bins HwsRomRcSensConfigHwsAndRadio                            = { [ (('h4000fc46 - 'h4000fc00) >> 1) : ((('h4000fc46 - 'h4000fc00 + 'd12) >> 1) - 1) ] };
    bins HwsRomRcSensActivation                                   = { [ (('h4000fc52 - 'h4000fc00) >> 1) : ((('h4000fc52 - 'h4000fc00 + 'd6) >> 1) - 1) ] };
    bins HwsRomRcSensPopulateOvlB2B                               = { [ (('h4000fc58 - 'h4000fc00) >> 1) : ((('h4000fc58 - 'h4000fc00 + 'd4) >> 1) - 1) ] };
    bins HwsRomCleActivationForFllOperation                       = { [ (('h4000fc5c - 'h4000fc00) >> 1) : ((('h4000fc5c - 'h4000fc00 + 'd14) >> 1) - 1) ] };
    bins HwsRomCleActivationForWkupOperation                      = { [ (('h4000fc6a - 'h4000fc00) >> 1) : ((('h4000fc6a - 'h4000fc00 + 'd14) >> 1) - 1) ] };
    bins HwsRomFsmDfMeasActivateB2B                               = { [ (('h4000fc78 - 'h4000fc00) >> 1) : ((('h4000fc78 - 'h4000fc00 + 'd16) >> 1) - 1) ] };
    bins HwsRomFsmFmuLoDivSymConfigHwsAndRadio                    = { [ (('h4000fc88 - 'h4000fc00) >> 1) : ((('h4000fc88 - 'h4000fc00 + 'd14) >> 1) - 1) ] };
    bins HwsRomFsmFmuLoDivSymVsSocActivateB2B                     = { [ (('h4000fc96 - 'h4000fc00) >> 1) : ((('h4000fc96 - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomEnvdetClkMeas                                      = { [ (('h4000fc9e - 'h4000fc00) >> 1) : ((('h4000fc9e - 'h4000fc00 + 'd12) >> 1) - 1) ] };
    bins HwsRomRtcClkMeas                                         = { [ (('h4000fcaa - 'h4000fc00) >> 1) : ((('h4000fcaa - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomSetAdbConfigForContWkup                            = { [ (('h4000fcb4 - 'h4000fc00) >> 1) : ((('h4000fcb4 - 'h4000fc00 + 'd6) >> 1) - 1) ] };
    bins HwsRomRestoreAdbConfigAfterContWkup                      = { [ (('h4000fcba - 'h4000fc00) >> 1) : ((('h4000fcba - 'h4000fc00 + 'd6) >> 1) - 1) ] };
    bins HwsRomPreAuxMeasSequence                                 = { [ (('h4000fcc0 - 'h4000fc00) >> 1) : ((('h4000fcc0 - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomPostAuxMeasSequence                                = { [ (('h4000fcc8 - 'h4000fc00) >> 1) : ((('h4000fcc8 - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomAuxMeasPopulateOvlB2B                              = { [ (('h4000fcd2 - 'h4000fc00) >> 1) : ((('h4000fcd2 - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomSymMeasPopulateOvlB2B                              = { [ (('h4000fcdc - 'h4000fc00) >> 1) : ((('h4000fcdc - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomFsmAuxMeasRxConfigClbAndRadio                      = { [ (('h4000fce4 - 'h4000fc00) >> 1) : ((('h4000fce4 - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomFsmAuxMeasRxConfigClbAndRadioForContWkup           = { [ (('h4000fcee - 'h4000fc00) >> 1) : ((('h4000fcee - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomFsmAuxMeasLoConfigClbAndRadio                      = { [ (('h4000fcf8 - 'h4000fc00) >> 1) : ((('h4000fcf8 - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomFsmSymMeasLoConfigClbAndRadio                      = { [ (('h4000fd02 - 'h4000fc00) >> 1) : ((('h4000fd02 - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomFsmSymMeasLcConfigClbAndRadio                      = { [ (('h4000fd0c - 'h4000fc00) >> 1) : ((('h4000fd0c - 'h4000fc00 + 'd14) >> 1) - 1) ] };
    bins HwsRomFsmMeasLoVrefVbpCalibConfigClbAndRadio             = { [ (('h4000fd1a - 'h4000fc00) >> 1) : ((('h4000fd1a - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomFsmMeasLoVrefVbpCalibConfigClbAndRadioNoSampling   = { [ (('h4000fd24 - 'h4000fc00) >> 1) : ((('h4000fd24 - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomFsmDfMeasConfigClbAndRadio                         = { [ (('h4000fd2e - 'h4000fc00) >> 1) : ((('h4000fd2e - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomFsmFllMeasActivateB2B                              = { [ (('h4000fd38 - 'h4000fc00) >> 1) : ((('h4000fd38 - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomFsmFllMeasActivateForContWkupB2B                   = { [ (('h4000fd40 - 'h4000fc00) >> 1) : ((('h4000fd40 - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomLoCalibPopulateOvlB2B                              = { [ (('h4000fd4a - 'h4000fc00) >> 1) : ((('h4000fd4a - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomFsmLoCalibConfigClbAndRadio                        = { [ (('h4000fd52 - 'h4000fc00) >> 1) : ((('h4000fd52 - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomFsmFllLoCalibActivateB2B                           = { [ (('h4000fd5c - 'h4000fc00) >> 1) : ((('h4000fd5c - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomFsmLoCalibLvNoOtp                                  = { [ (('h4000fd64 - 'h4000fc00) >> 1) : ((('h4000fd64 - 'h4000fc00 + 'd18) >> 1) - 1) ] };
    bins HwsRomSymCalibPopulateOvlB2B                             = { [ (('h4000fd76 - 'h4000fc00) >> 1) : ((('h4000fd76 - 'h4000fc00 + 'd6) >> 1) - 1) ] };
    bins HwsRomFsmSymCalibConfigClbAndRadio                       = { [ (('h4000fd7c - 'h4000fc00) >> 1) : ((('h4000fd7c - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomFsmFllSymCalibActivateB2B                          = { [ (('h4000fd86 - 'h4000fc00) >> 1) : ((('h4000fd86 - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomEncryptDataB2B                                     = { [ (('h4000fd8e - 'h4000fc00) >> 1) : ((('h4000fd8e - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomFsmPgxConfigHwsAndRadio                            = { [ (('h4000fd98 - 'h4000fc00) >> 1) : ((('h4000fd98 - 'h4000fc00 + 'd12) >> 1) - 1) ] };
    bins HwsRomFsmPgxLoDivSymConfigHwsAndRadio                    = { [ (('h4000fda4 - 'h4000fc00) >> 1) : ((('h4000fda4 - 'h4000fc00 + 'd14) >> 1) - 1) ] };
    bins HwsRomFsmPgxLoDivSymForBle5ConfigHwsAndRadio             = { [ (('h4000fdb2 - 'h4000fc00) >> 1) : ((('h4000fdb2 - 'h4000fc00 + 'd20) >> 1) - 1) ] };
    bins HwsRomFsmPgxActivateMfgId                                = { [ (('h4000fdc6 - 'h4000fc00) >> 1) : ((('h4000fdc6 - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomFsmPgxActivateSrvcId                               = { [ (('h4000fdce - 'h4000fc00) >> 1) : ((('h4000fdce - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomFsmPgxActivateRawNonWhiteLegacy                    = { [ (('h4000fdd6 - 'h4000fc00) >> 1) : ((('h4000fdd6 - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomFsmPgxActivateAdvExtInd                            = { [ (('h4000fdde - 'h4000fc00) >> 1) : ((('h4000fdde - 'h4000fc00 + 'd10) >> 1) - 1) ] };
    bins HwsRomFsmPgxActivateAdvExtIndB2B                         = { [ (('h4000fde8 - 'h4000fc00) >> 1) : ((('h4000fde8 - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomFsmPgxActivateAuxAdvInd                            = { [ (('h4000fdf0 - 'h4000fc00) >> 1) : ((('h4000fdf0 - 'h4000fc00 + 'd16) >> 1) - 1) ] };
    bins HwsRomFsmPgxActivateAuxAdvIndRaw                         = { [ (('h4000fe00 - 'h4000fc00) >> 1) : ((('h4000fe00 - 'h4000fc00 + 'd18) >> 1) - 1) ] };
    bins HwsRomFsmPgxActivateMfgIdNoOtp                           = { [ (('h4000fe12 - 'h4000fc00) >> 1) : ((('h4000fe12 - 'h4000fc00 + 'd18) >> 1) - 1) ] };
    bins HwsRomFsmPgxActivateSrvcIdNoOtp                          = { [ (('h4000fe24 - 'h4000fc00) >> 1) : ((('h4000fe24 - 'h4000fc00 + 'd18) >> 1) - 1) ] };
    bins HwsRomPreparePacketWithConstsB2B                         = { [ (('h4000fe36 - 'h4000fc00) >> 1) : ((('h4000fe36 - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomRadioTrngB2B                                       = { [ (('h4000fe3e - 'h4000fc00) >> 1) : ((('h4000fe3e - 'h4000fc00 + 'd20) >> 1) - 1) ] };
    bins HwsRomRetWkupWithFreqOffset                              = { [ (('h4000fe52 - 'h4000fc00) >> 1) : ((('h4000fe52 - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomContWkupWithFreqOffset                             = { [ (('h4000fe5a - 'h4000fc00) >> 1) : ((('h4000fe5a - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomRetWkupWithFreqOffsetWithException                 = { [ (('h4000fe62 - 'h4000fc00) >> 1) : ((('h4000fe62 - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomContWkupWithFreqOffsetWithException                = { [ (('h4000fe6a - 'h4000fc00) >> 1) : ((('h4000fe6a - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins HwsRomLoProxSensingInit                                  = { [ (('h4000fe72 - 'h4000fc00) >> 1) : ((('h4000fe72 - 'h4000fc00 + 'd14) >> 1) - 1) ] };
    bins HwsRomLoProxSensingExecute                               = { [ (('h4000fe80 - 'h4000fc00) >> 1) : ((('h4000fe80 - 'h4000fc00 + 'd20) >> 1) - 1) ] };
    bins HwsRomSymCalib                                           = { [ (('h4000fe94 - 'h4000fc00) >> 1) : ((('h4000fe94 - 'h4000fc00 + 'd26) >> 1) - 1) ] };
    bins HwsRomPowerGearing                                       = { [ (('h4000feae - 'h4000fc00) >> 1) : ((('h4000feae - 'h4000fc00 + 'd24) >> 1) - 1) ] };
    bins PowerGearingExit                                         = { [ (('h4000fec2 - 'h4000fc00) >> 1) : ((('h4000fec2 - 'h4000fc00 + 'd20) >> 1) - 1) ] };
    bins HwsRomLcAuxIdacCalibInit                                 = { [ (('h4000fec6 - 'h4000fc00) >> 1) : ((('h4000fec6 - 'h4000fc00 + 'd12) >> 1) - 1) ] };
    bins HwsRomLcAuxIdacCalibExecute                              = { [ (('h4000fed2 - 'h4000fc00) >> 1) : ((('h4000fed2 - 'h4000fc00 + 'd36) >> 1) - 1) ] };
    bins LcAuxIdacCalibExecute                                    = { [ (('h4000fed2 - 'h4000fc00) >> 1) : ((('h4000fed2 - 'h4000fc00 + 'd0) >> 1) - 1) ] };
    bins HwsRomPreHarvesterFlow                                   = { [ (('h4000fef6 - 'h4000fc00) >> 1) : ((('h4000fef6 - 'h4000fc00 + 'd8) >> 1) - 1) ] };
    bins RAW_TX_LOOP                                              = { [ (('h4000fefe - 'h4000fc00) >> 1) : ((('h4000fefe - 'h4000fc00 + 'd44) >> 1) - 1) ] };
    bins repeat_tx_loop                                           = { [ (('h4000ff0e - 'h4000fc00) >> 1) : ((('h4000ff0e - 'h4000fc00 + 'd16) >> 1) - 1) ] };
    bins HarvesterTxStart                                         = { [ (('h4000ff22 - 'h4000fc00) >> 1) : ((('h4000ff22 - 'h4000fc00 + 'd36) >> 1) - 1) ] };
    bins EndHarvFlow                                              = { [ (('h4000ff28 - 'h4000fc00) >> 1) : ((('h4000ff28 - 'h4000fc00 + 'd42) >> 1) - 1) ] };
    bins FlowManagerFsm                                           = { [ (('h40010e0c - 'h4000fc00) >> 1) : ((('h40010e0c - 'h4000fc00 + 'd12) >> 1) - 1) ] };
    bins TempSensingLoop                                          = { [ (('h40010e3c - 'h4000fc00) >> 1) : ((('h40010e3c - 'h4000fc00 + 'd60) >> 1) - 1) ] };
    bins TempSensingLoopExecute                                   = { [ (('h40010e42 - 'h4000fc00) >> 1) : ((('h40010e42 - 'h4000fc00 + 'd66) >> 1) - 1) ] };
    bins LoProxSensingLoop                                        = { [ (('h40010e4c - 'h4000fc00) >> 1) : ((('h40010e4c - 'h4000fc00 + 'd76) >> 1) - 1) ] };
    bins RcSensorLoop                                             = { [ (('h40010e52 - 'h4000fc00) >> 1) : ((('h40010e52 - 'h4000fc00 + 'd82) >> 1) - 1) ] };
    bins RcSensorLoopExecute                                      = { [ (('h40010e5a - 'h4000fc00) >> 1) : ((('h40010e5a - 'h4000fc00 + 'd90) >> 1) - 1) ] };
    bins TamperSensingLoop                                        = { [ (('h40010e64 - 'h4000fc00) >> 1) : ((('h40010e64 - 'h4000fc00 + 'd100) >> 1) - 1) ] };
    bins SystemClksMeasLoop                                       = { [ (('h40010e6a - 'h4000fc00) >> 1) : ((('h40010e6a - 'h4000fc00 + 'd106) >> 1) - 1) ] };
    bins SystemClksMeasExecute                                    = { [ (('h40010e6e - 'h4000fc00) >> 1) : ((('h40010e6e - 'h4000fc00 + 'd110) >> 1) - 1) ] };
    bins SocMeasLoop                                              = { [ (('h40010e76 - 'h4000fc00) >> 1) : ((('h40010e76 - 'h4000fc00 + 'd118) >> 1) - 1) ] };
    bins EnvdetMeasLoop                                           = { [ (('h40010e7e - 'h4000fc00) >> 1) : ((('h40010e7e - 'h4000fc00 + 'd126) >> 1) - 1) ] };
    bins RtcMeasLoop                                              = { [ (('h40010e86 - 'h4000fc00) >> 1) : ((('h40010e86 - 'h4000fc00 + 'd134) >> 1) - 1) ] };
    bins RxSweepAndAuxMeasLoop                                    = { [ (('h40010e90 - 'h4000fc00) >> 1) : ((('h40010e90 - 'h4000fc00 + 'd144) >> 1) - 1) ] };
    bins RxSweep                                                  = { [ (('h40010e9a - 'h4000fc00) >> 1) : ((('h40010e9a - 'h4000fc00 + 'd154) >> 1) - 1) ] };
    bins AuxMeas                                                  = { [ (('h40010ea4 - 'h4000fc00) >> 1) : ((('h40010ea4 - 'h4000fc00 + 'd164) >> 1) - 1) ] };
    bins AuxMeasExecute                                           = { [ (('h40010eae - 'h4000fc00) >> 1) : ((('h40010eae - 'h4000fc00 + 'd174) >> 1) - 1) ] };
    bins PostAuxMeas                                              = { [ (('h40010eb6 - 'h4000fc00) >> 1) : ((('h40010eb6 - 'h4000fc00 + 'd182) >> 1) - 1) ] };
    bins PostRxSweepAndAuxMeas                                    = { [ (('h40010eb8 - 'h4000fc00) >> 1) : ((('h40010eb8 - 'h4000fc00 + 'd184) >> 1) - 1) ] };
    bins LoTxRxCalibLoop                                          = { [ (('h40010ebc - 'h4000fc00) >> 1) : ((('h40010ebc - 'h4000fc00 + 'd188) >> 1) - 1) ] };
    bins LoTxRxCalibExecute                                       = { [ (('h40010ec2 - 'h4000fc00) >> 1) : ((('h40010ec2 - 'h4000fc00 + 'd194) >> 1) - 1) ] };
    bins SymCalibLoop                                             = { [ (('h40010ece - 'h4000fc00) >> 1) : ((('h40010ece - 'h4000fc00 + 'd206) >> 1) - 1) ] };
    bins SecAndTxLoop                                             = { [ (('h40010ed2 - 'h4000fc00) >> 1) : ((('h40010ed2 - 'h4000fc00 + 'd210) >> 1) - 1) ] };
    bins TxSprinkler                                              = { [ (('h40010edc - 'h4000fc00) >> 1) : ((('h40010edc - 'h4000fc00 + 'd220) >> 1) - 1) ] };
    bins PreparePacketLoop                                        = { [ (('h40010ee4 - 'h4000fc00) >> 1) : ((('h40010ee4 - 'h4000fc00 + 'd228) >> 1) - 1) ] };
    bins TxLegacyLoop                                             = { [ (('h40010ef4 - 'h4000fc00) >> 1) : ((('h40010ef4 - 'h4000fc00 + 'd244) >> 1) - 1) ] };
    bins TxBle5Loop                                               = { [ (('h40010f02 - 'h4000fc00) >> 1) : ((('h40010f02 - 'h4000fc00 + 'd258) >> 1) - 1) ] };
    bins TempStaticCompLoop                                       = { [ (('h40010f1a - 'h4000fc00) >> 1) : ((('h40010f1a - 'h4000fc00 + 'd282) >> 1) - 1) ] };
    bins PowerGearingLoop                                         = { [ (('h40010f20 - 'h4000fc00) >> 1) : ((('h40010f20 - 'h4000fc00 + 'd288) >> 1) - 1) ] };
    bins LcAuxIdacCalibLoop                                       = { [ (('h40010f24 - 'h4000fc00) >> 1) : ((('h40010f24 - 'h4000fc00 + 'd292) >> 1) - 1) ] };
    bins WkupThresholdCalibLoop                                   = { [ (('h40010f2a - 'h4000fc00) >> 1) : ((('h40010f2a - 'h4000fc00 + 'd298) >> 1) - 1) ] };
    bins WkupLowSensitivityCalib                                  = { [ (('h40010f30 - 'h4000fc00) >> 1) : ((('h40010f30 - 'h4000fc00 + 'd304) >> 1) - 1) ] };
    bins LoVrefVbpCalibLoop                                       = { [ (('h40010f3a - 'h4000fc00) >> 1) : ((('h40010f3a - 'h4000fc00 + 'd314) >> 1) - 1) ] };
    bins LoVrefVbpCalibExecute                                    = { [ (('h40010f40 - 'h4000fc00) >> 1) : ((('h40010f40 - 'h4000fc00 + 'd320) >> 1) - 1) ] };
    bins ModIdxCalibLoop                                          = { [ (('h40010f4e - 'h4000fc00) >> 1) : ((('h40010f4e - 'h4000fc00 + 'd334) >> 1) - 1) ] };
    bins ModIdxCalibExecute                                       = { [ (('h40010f54 - 'h4000fc00) >> 1) : ((('h40010f54 - 'h4000fc00 + 'd340) >> 1) - 1) ] };
    bins MiniRxLoop                                               = { [ (('h40010f60 - 'h4000fc00) >> 1) : ((('h40010f60 - 'h4000fc00 + 'd352) >> 1) - 1) ] };
    bins MiniRxMainLoop                                           = { [ (('h40010f6c - 'h4000fc00) >> 1) : ((('h40010f6c - 'h4000fc00 + 'd364) >> 1) - 1) ] };
    bins NoContWuForFirstRun                                      = { [ (('h40010f6e - 'h4000fc00) >> 1) : ((('h40010f6e - 'h4000fc00 + 'd366) >> 1) - 1) ] };
    bins ExitCheckRx                                              = { [ (('h40010f7e - 'h4000fc00) >> 1) : ((('h40010f7e - 'h4000fc00 + 'd382) >> 1) - 1) ] };
    bins HarvesterFlow                                            = { [ (('h40010f88 - 'h4000fc00) >> 1) : ((('h40010f88 - 'h4000fc00 + 'd392) >> 1) - 1) ] };