    bins SpuRomRadioModeForTxLv                           = { [ (('h4000d668 - 'h4000d668) >> 1) : ((('h4000d668 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForTxLv                           = { [ (('h4000d670 - 'h4000d668) >> 1) : ((('h4000d670 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForTxHv                           = { [ (('h4000d688 - 'h4000d668) >> 1) : ((('h4000d688 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForTxHv                           = { [ (('h4000d690 - 'h4000d668) >> 1) : ((('h4000d690 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForSymCalibLv                     = { [ (('h4000d6a8 - 'h4000d668) >> 1) : ((('h4000d6a8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForSymCalibLv                     = { [ (('h4000d6b0 - 'h4000d668) >> 1) : ((('h4000d6b0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForSymCalibHv                     = { [ (('h4000d6c8 - 'h4000d668) >> 1) : ((('h4000d6c8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForSymCalibHv                     = { [ (('h4000d6d0 - 'h4000d668) >> 1) : ((('h4000d6d0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForLoCalibLv                      = { [ (('h4000d6e8 - 'h4000d668) >> 1) : ((('h4000d6e8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForLoCalibLv                      = { [ (('h4000d6f0 - 'h4000d668) >> 1) : ((('h4000d6f0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForLoCalibHv                      = { [ (('h4000d708 - 'h4000d668) >> 1) : ((('h4000d708 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForLoCalibHv                      = { [ (('h4000d710 - 'h4000d668) >> 1) : ((('h4000d710 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForMeasureLv                      = { [ (('h4000d728 - 'h4000d668) >> 1) : ((('h4000d728 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForMeasureLv                      = { [ (('h4000d730 - 'h4000d668) >> 1) : ((('h4000d730 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForMeasureHv                      = { [ (('h4000d748 - 'h4000d668) >> 1) : ((('h4000d748 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForMeasureHv                      = { [ (('h4000d750 - 'h4000d668) >> 1) : ((('h4000d750 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForMeasureLC                      = { [ (('h4000d768 - 'h4000d668) >> 1) : ((('h4000d768 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForMeasureLC                      = { [ (('h4000d770 - 'h4000d668) >> 1) : ((('h4000d770 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForTempSensLv                     = { [ (('h4000d788 - 'h4000d668) >> 1) : ((('h4000d788 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForTempSensLv                     = { [ (('h4000d790 - 'h4000d668) >> 1) : ((('h4000d790 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForRcSensCap                      = { [ (('h4000d7a8 - 'h4000d668) >> 1) : ((('h4000d7a8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForRcSensCap                      = { [ (('h4000d7b0 - 'h4000d668) >> 1) : ((('h4000d7b0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForRcSensRes                      = { [ (('h4000d7c8 - 'h4000d668) >> 1) : ((('h4000d7c8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForRcSensRes                      = { [ (('h4000d7d0 - 'h4000d668) >> 1) : ((('h4000d7d0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForLoDivSymLv                     = { [ (('h4000d7e8 - 'h4000d668) >> 1) : ((('h4000d7e8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForLoDivSymLv                     = { [ (('h4000d7f0 - 'h4000d668) >> 1) : ((('h4000d7f0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForLoDivSymHv                     = { [ (('h4000d808 - 'h4000d668) >> 1) : ((('h4000d808 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForLoDivSymHv                     = { [ (('h4000d810 - 'h4000d668) >> 1) : ((('h4000d810 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForLoVrefVbpCalibLv               = { [ (('h4000d828 - 'h4000d668) >> 1) : ((('h4000d828 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForLoVrefVbpCalibLv               = { [ (('h4000d830 - 'h4000d668) >> 1) : ((('h4000d830 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForLoVrefVbpCalibHv               = { [ (('h4000d848 - 'h4000d668) >> 1) : ((('h4000d848 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForLoVrefVbpCalibHv               = { [ (('h4000d850 - 'h4000d668) >> 1) : ((('h4000d850 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForTxlvDFmeas                     = { [ (('h4000d868 - 'h4000d668) >> 1) : ((('h4000d868 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForTxlvDFmeas                     = { [ (('h4000d870 - 'h4000d668) >> 1) : ((('h4000d870 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForTxhvDFmeas                     = { [ (('h4000d888 - 'h4000d668) >> 1) : ((('h4000d888 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForTxhvDFmeas                     = { [ (('h4000d890 - 'h4000d668) >> 1) : ((('h4000d890 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioModeForRng_lo                         = { [ (('h4000d8a8 - 'h4000d668) >> 1) : ((('h4000d8a8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioInitForRng_lo                         = { [ (('h4000d8b0 - 'h4000d668) >> 1) : ((('h4000d8b0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomMemCopyRadioInit                           = { [ (('h4000d8c8 - 'h4000d668) >> 1) : ((('h4000d8c8 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomRadioInit                                  = { [ (('h4000d8e0 - 'h4000d668) >> 1) : ((('h4000d8e0 - 'h4000d668 + 'd40) >> 1) - 1) ] };
    bins SpuRomHwsLinkPreJump                             = { [ (('h4000d908 - 'h4000d668) >> 1) : ((('h4000d908 - 'h4000d668 + 'd48) >> 1) - 1) ] };
    bins SpuRomHwsLinkPostJump                            = { [ (('h4000d938 - 'h4000d668) >> 1) : ((('h4000d938 - 'h4000d668 + 'd52) >> 1) - 1) ] };
    bins SpuRomExceptionHandler                           = { [ (('h4000d970 - 'h4000d668) >> 1) : ((('h4000d970 - 'h4000d668 + 'd128) >> 1) - 1) ] };
    bins SpuRomJumpXRdrsFromNet                           = { [ (('h4000d9f0 - 'h4000d668) >> 1) : ((('h4000d9f0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomJumpXRdrsRelativeToEndFromNet              = { [ (('h4000da08 - 'h4000d668) >> 1) : ((('h4000da08 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomJumpXRdrsFromRrt                           = { [ (('h4000da20 - 'h4000d668) >> 1) : ((('h4000da20 - 'h4000d668 + 'd40) >> 1) - 1) ] };
    bins SpuRomJumpXRdrsRelativeToEndFromRrt              = { [ (('h4000da48 - 'h4000d668) >> 1) : ((('h4000da48 - 'h4000d668 + 'd36) >> 1) - 1) ] };
    bins SpuRomHwsJumpToSpecificRdr                       = { [ (('h4000da70 - 'h4000d668) >> 1) : ((('h4000da70 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomJumpXRdrs                                  = { [ (('h4000da88 - 'h4000d668) >> 1) : ((('h4000da88 - 'h4000d668 + 'd16) >> 1) - 1) ] };
    bins SpuRomJumpXRdrsRelativeToEnd                     = { [ (('h4000da98 - 'h4000d668) >> 1) : ((('h4000da98 - 'h4000d668 + 'd16) >> 1) - 1) ] };
    bins SpuRomSecCopyKeysFromOtp                         = { [ (('h4000daa8 - 'h4000d668) >> 1) : ((('h4000daa8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SPU_SecDMAPreFetch                               = { [ (('h4000dab0 - 'h4000d668) >> 1) : ((('h4000dab0 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomSecPreFetch                                = { [ (('h4000dac0 - 'h4000d668) >> 1) : ((('h4000dac0 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SPU_SecProcess                                   = { [ (('h4000dad0 - 'h4000d668) >> 1) : ((('h4000dad0 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SPU_SecDMAPush                                   = { [ (('h4000dae0 - 'h4000d668) >> 1) : ((('h4000dae0 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomSecPush                                    = { [ (('h4000dae8 - 'h4000d668) >> 1) : ((('h4000dae8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomInitFromGnvm                               = { [ (('h4000daf0 - 'h4000d668) >> 1) : ((('h4000daf0 - 'h4000d668 + 'd64) >> 1) - 1) ] };
    bins SpuRomClearIspExcpFlags                          = { [ (('h4000db30 - 'h4000d668) >> 1) : ((('h4000db30 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomDummy                                      = { [ (('h4000db48 - 'h4000d668) >> 1) : ((('h4000db48 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomDontIncTOctrInExcp                         = { [ (('h4000db50 - 'h4000d668) >> 1) : ((('h4000db50 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomIncTOctrInExcp                             = { [ (('h4000db58 - 'h4000d668) >> 1) : ((('h4000db58 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomSetStateOperationDoneInd                   = { [ (('h4000db60 - 'h4000d668) >> 1) : ((('h4000db60 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomClearStateOperationDoneInd                 = { [ (('h4000db68 - 'h4000d668) >> 1) : ((('h4000db68 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins Spu_TempSensorSrrInit                            = { [ (('h4000db70 - 'h4000d668) >> 1) : ((('h4000db70 - 'h4000d668 + 'd160) >> 1) - 1) ] };
    bins Spu_TempSensor_dig_ctl_srr                       = { [ (('h4000dc10 - 'h4000d668) >> 1) : ((('h4000dc10 - 'h4000d668 + 'd212) >> 1) - 1) ] };
    bins Spu_TempSensorInit                               = { [ (('h4000dce8 - 'h4000d668) >> 1) : ((('h4000dce8 - 'h4000d668 + 'd116) >> 1) - 1) ] };
    bins Spu_TempSensor_dig_ctl                           = { [ (('h4000dd60 - 'h4000d668) >> 1) : ((('h4000dd60 - 'h4000d668 + 'd184) >> 1) - 1) ] };
    bins Spu_TempSensor_analog_ctl                        = { [ (('h4000de18 - 'h4000d668) >> 1) : ((('h4000de18 - 'h4000d668 + 'd204) >> 1) - 1) ] };
    bins Spu_TempSensor_first_boot_ctl                    = { [ (('h4000dee8 - 'h4000d668) >> 1) : ((('h4000dee8 - 'h4000d668 + 'd44) >> 1) - 1) ] };
    bins Spu_TempSensor_ctl                               = { [ (('h4000df18 - 'h4000d668) >> 1) : ((('h4000df18 - 'h4000d668 + 'd48) >> 1) - 1) ] };
    bins Spu_TempSensorInit_ctl                           = { [ (('h4000df48 - 'h4000d668) >> 1) : ((('h4000df48 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomConfigClbForTempSense                      = { [ (('h4000df60 - 'h4000d668) >> 1) : ((('h4000df60 - 'h4000d668 + 'd44) >> 1) - 1) ] };
    bins SpuRomTempSensorCfgOtpToOvl                      = { [ (('h4000df90 - 'h4000d668) >> 1) : ((('h4000df90 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRcSensCfgOtpToOvl                          = { [ (('h4000df98 - 'h4000d668) >> 1) : ((('h4000df98 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomConfigHwsForRcSensing                      = { [ (('h4000dfa0 - 'h4000d668) >> 1) : ((('h4000dfa0 - 'h4000d668 + 'd48) >> 1) - 1) ] };
    bins SpuRomRcSensSetParams                            = { [ (('h4000dfd0 - 'h4000d668) >> 1) : ((('h4000dfd0 - 'h4000d668 + 'd36) >> 1) - 1) ] };
    bins SpuRomRcMaskLc                                   = { [ (('h4000dff8 - 'h4000d668) >> 1) : ((('h4000dff8 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRcSensFunc                                 = { [ (('h4000e010 - 'h4000d668) >> 1) : ((('h4000e010 - 'h4000d668 + 'd36) >> 1) - 1) ] };
    bins SpuRomDisableRadioTurnOff                        = { [ (('h4000e038 - 'h4000d668) >> 1) : ((('h4000e038 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomEnableRadioTurnOff                         = { [ (('h4000e040 - 'h4000d668) >> 1) : ((('h4000e040 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomSetRadioForTx                              = { [ (('h4000e048 - 'h4000d668) >> 1) : ((('h4000e048 - 'h4000d668 + 'd52) >> 1) - 1) ] };
    bins SpuRomSetRadioForSymCalib                        = { [ (('h4000e080 - 'h4000d668) >> 1) : ((('h4000e080 - 'h4000d668 + 'd52) >> 1) - 1) ] };
    bins SpuRomSetRadioForLoCalib                         = { [ (('h4000e0b8 - 'h4000d668) >> 1) : ((('h4000e0b8 - 'h4000d668 + 'd52) >> 1) - 1) ] };
    bins SpuRomSetRadioForMeasure                         = { [ (('h4000e0f0 - 'h4000d668) >> 1) : ((('h4000e0f0 - 'h4000d668 + 'd52) >> 1) - 1) ] };
    bins SpuRomSetRadioForRcSens                          = { [ (('h4000e128 - 'h4000d668) >> 1) : ((('h4000e128 - 'h4000d668 + 'd52) >> 1) - 1) ] };
    bins SpuRomSetRadioForLoDivSym                        = { [ (('h4000e160 - 'h4000d668) >> 1) : ((('h4000e160 - 'h4000d668 + 'd52) >> 1) - 1) ] };
    bins SpuRomSetRadioForMeasLoVrefVbpCalib              = { [ (('h4000e198 - 'h4000d668) >> 1) : ((('h4000e198 - 'h4000d668 + 'd28) >> 1) - 1) ] };
    bins SpuRomSetRadioForMeasLoVrefVbpCalibNoSampling    = { [ (('h4000e1b8 - 'h4000d668) >> 1) : ((('h4000e1b8 - 'h4000d668 + 'd52) >> 1) - 1) ] };
    bins SpuRomSetRadioForDFmeas                          = { [ (('h4000e1f0 - 'h4000d668) >> 1) : ((('h4000e1f0 - 'h4000d668 + 'd52) >> 1) - 1) ] };
    bins SpuRomTurnOtpPowerOn                             = { [ (('h4000e228 - 'h4000d668) >> 1) : ((('h4000e228 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomTurnOtpPowerOff                            = { [ (('h4000e230 - 'h4000d668) >> 1) : ((('h4000e230 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomReduceSramAndRomDcdcFreq                   = { [ (('h4000e238 - 'h4000d668) >> 1) : ((('h4000e238 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomSetActiveClkDividerRatioToMax              = { [ (('h4000e248 - 'h4000d668) >> 1) : ((('h4000e248 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomRestoreActiveClkDividerRatio               = { [ (('h4000e258 - 'h4000d668) >> 1) : ((('h4000e258 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins Populate_Radio_ISP                               = { [ (('h4000e270 - 'h4000d668) >> 1) : ((('h4000e270 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins Populate_Radio_HWS                               = { [ (('h4000e278 - 'h4000d668) >> 1) : ((('h4000e278 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins Copy_AuxMeas_OTP_To_scratch                      = { [ (('h4000e280 - 'h4000d668) >> 1) : ((('h4000e280 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SPU_SET_Measurement_Configuration                = { [ (('h4000e288 - 'h4000d668) >> 1) : ((('h4000e288 - 'h4000d668 + 'd28) >> 1) - 1) ] };
    bins Copy_LoCalib_OTP_To_scratch                      = { [ (('h4000e2a8 - 'h4000d668) >> 1) : ((('h4000e2a8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SPU_SET_LO_Calibration_Configuration             = { [ (('h4000e2b0 - 'h4000d668) >> 1) : ((('h4000e2b0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins Copy_SymCalib_OTP_To_scratch                     = { [ (('h4000e2c8 - 'h4000d668) >> 1) : ((('h4000e2c8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SPU_SET_Sym_Calibration_Configuration            = { [ (('h4000e2d0 - 'h4000d668) >> 1) : ((('h4000e2d0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SPU_SET_PGX_Configuration                        = { [ (('h4000e2e8 - 'h4000d668) >> 1) : ((('h4000e2e8 - 'h4000d668 + 'd32) >> 1) - 1) ] };
    bins Copy_Measurement_To_ISP                          = { [ (('h4000e308 - 'h4000d668) >> 1) : ((('h4000e308 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins Copy_DataKeys_OTP_To_scratch                     = { [ (('h4000e310 - 'h4000d668) >> 1) : ((('h4000e310 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins Copy_IDKeys_OTP_To_scratch                       = { [ (('h4000e318 - 'h4000d668) >> 1) : ((('h4000e318 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SPU_CopyTRNGToISP                                = { [ (('h4000e320 - 'h4000d668) >> 1) : ((('h4000e320 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SPU_PopulatePGX                                  = { [ (('h4000e328 - 'h4000d668) >> 1) : ((('h4000e328 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomCloseWkup                                  = { [ (('h4000e330 - 'h4000d668) >> 1) : ((('h4000e330 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomSetWkupMode3                               = { [ (('h4000e348 - 'h4000d668) >> 1) : ((('h4000e348 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SPU_SetCCA                                       = { [ (('h4000e350 - 'h4000d668) >> 1) : ((('h4000e350 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomInitSwspad0To31                            = { [ (('h4000e360 - 'h4000d668) >> 1) : ((('h4000e360 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomInitSwspadGnvm                             = { [ (('h4000e378 - 'h4000d668) >> 1) : ((('h4000e378 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomInitSrr                                    = { [ (('h4000e380 - 'h4000d668) >> 1) : ((('h4000e380 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomInitHrr                                    = { [ (('h4000e398 - 'h4000d668) >> 1) : ((('h4000e398 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomCopyFrequentHrrGnvmToSrrOvl                = { [ (('h4000e3b0 - 'h4000d668) >> 1) : ((('h4000e3b0 - 'h4000d668 + 'd252) >> 1) - 1) ] };
    bins SpuRomCopyFrequentSwGnvmToSrrOvl                 = { [ (('h4000e4b0 - 'h4000d668) >> 1) : ((('h4000e4b0 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomInitAuxMeas                                = { [ (('h4000e4b8 - 'h4000d668) >> 1) : ((('h4000e4b8 - 'h4000d668 + 'd16) >> 1) - 1) ] };
    bins SpuRomInitClbContext0                            = { [ (('h4000e4c8 - 'h4000d668) >> 1) : ((('h4000e4c8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomInitClbSkipN                               = { [ (('h4000e4d0 - 'h4000d668) >> 1) : ((('h4000e4d0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomSetInitialParamsUntilFirstTempCompPart1    = { [ (('h4000e4e8 - 'h4000d668) >> 1) : ((('h4000e4e8 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomSetInitialParamsUntilFirstTempCompPart2    = { [ (('h4000e4f8 - 'h4000d668) >> 1) : ((('h4000e4f8 - 'h4000d668 + 'd68) >> 1) - 1) ] };
    bins SpuRomFirstBootInitUntilFirstTempComp            = { [ (('h4000e540 - 'h4000d668) >> 1) : ((('h4000e540 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRadioOtpToSrr                              = { [ (('h4000e558 - 'h4000d668) >> 1) : ((('h4000e558 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomRadioSrrToHws                              = { [ (('h4000e560 - 'h4000d668) >> 1) : ((('h4000e560 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomPgxOtpToSrr                                = { [ (('h4000e568 - 'h4000d668) >> 1) : ((('h4000e568 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomPgxSrrToHws                                = { [ (('h4000e570 - 'h4000d668) >> 1) : ((('h4000e570 - 'h4000d668 + 'd28) >> 1) - 1) ] };
    bins SpuRomPgxSrrToHws64Bit                           = { [ (('h4000e590 - 'h4000d668) >> 1) : ((('h4000e590 - 'h4000d668 + 'd52) >> 1) - 1) ] };
    bins SpuRomPgxSrrToHwsRaw128Bit                       = { [ (('h4000e5c8 - 'h4000d668) >> 1) : ((('h4000e5c8 - 'h4000d668 + 'd80) >> 1) - 1) ] };
    bins SpuRomPgxHwsToSrr                                = { [ (('h4000e618 - 'h4000d668) >> 1) : ((('h4000e618 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomSetRawPacketSize                           = { [ (('h4000e620 - 'h4000d668) >> 1) : ((('h4000e620 - 'h4000d668 + 'd28) >> 1) - 1) ] };
    bins SpuRomCopyRawPcktCrc                             = { [ (('h4000e640 - 'h4000d668) >> 1) : ((('h4000e640 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomCopyLoDivSymFromOvlToHws                   = { [ (('h4000e648 - 'h4000d668) >> 1) : ((('h4000e648 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomSetLoDivSymFromCh37InOvl                   = { [ (('h4000e650 - 'h4000d668) >> 1) : ((('h4000e650 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomSetLoDivSymFromCh37InClb                   = { [ (('h4000e658 - 'h4000d668) >> 1) : ((('h4000e658 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomSetAwdtSoftRguMaxTh                        = { [ (('h4000e660 - 'h4000d668) >> 1) : ((('h4000e660 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomTxBle5LengthJump                           = { [ (('h4000e678 - 'h4000d668) >> 1) : ((('h4000e678 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomSyncEnvDetWithSoc                          = { [ (('h4000e690 - 'h4000d668) >> 1) : ((('h4000e690 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomCopySrrToAuxPgxData                        = { [ (('h4000e698 - 'h4000d668) >> 1) : ((('h4000e698 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomSetWhtnForBle5                             = { [ (('h4000e6a0 - 'h4000d668) >> 1) : ((('h4000e6a0 - 'h4000d668 + 'd16) >> 1) - 1) ] };
    bins SpuRomSetPreambleAndDfSizeForBle5                = { [ (('h4000e6b0 - 'h4000d668) >> 1) : ((('h4000e6b0 - 'h4000d668 + 'd64) >> 1) - 1) ] };
    bins SpuRomSetPsuRadioClkDivForTx                     = { [ (('h4000e6f0 - 'h4000d668) >> 1) : ((('h4000e6f0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomRestorePsuRadioClkDivAfterTx               = { [ (('h4000e708 - 'h4000d668) >> 1) : ((('h4000e708 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomHwsOtpToHrr                                = { [ (('h4000e720 - 'h4000d668) >> 1) : ((('h4000e720 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomAuxMeasOtpToIsp                            = { [ (('h4000e730 - 'h4000d668) >> 1) : ((('h4000e730 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomAuxMeasIspToOvl                            = { [ (('h4000e738 - 'h4000d668) >> 1) : ((('h4000e738 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomAuxMeasMsrCtl12ToOvl                       = { [ (('h4000e740 - 'h4000d668) >> 1) : ((('h4000e740 - 'h4000d668 + 'd16) >> 1) - 1) ] };
    bins SpuRomSymMeasMsrCtl12ToOvl                       = { [ (('h4000e750 - 'h4000d668) >> 1) : ((('h4000e750 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomAuxMeasResOvlToIsp                         = { [ (('h4000e768 - 'h4000d668) >> 1) : ((('h4000e768 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomAuxMeasResIspToOvl                         = { [ (('h4000e770 - 'h4000d668) >> 1) : ((('h4000e770 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomAuxMeasResOvlToClb                         = { [ (('h4000e778 - 'h4000d668) >> 1) : ((('h4000e778 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomClbContextOtpToSrr                         = { [ (('h4000e780 - 'h4000d668) >> 1) : ((('h4000e780 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomClbContextSrrToOvl                         = { [ (('h4000e790 - 'h4000d668) >> 1) : ((('h4000e790 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomClbContextOvlToClb                         = { [ (('h4000e7a0 - 'h4000d668) >> 1) : ((('h4000e7a0 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomAuxMeasCfgOtpToOvl                         = { [ (('h4000e7a8 - 'h4000d668) >> 1) : ((('h4000e7a8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomAuxMeasOvlToClb                            = { [ (('h4000e7b0 - 'h4000d668) >> 1) : ((('h4000e7b0 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomLoCalibOtpToOvl                            = { [ (('h4000e7b8 - 'h4000d668) >> 1) : ((('h4000e7b8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomLoCalibOvlToClb                            = { [ (('h4000e7c0 - 'h4000d668) >> 1) : ((('h4000e7c0 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomSymCalibOtpToOvl                           = { [ (('h4000e7c8 - 'h4000d668) >> 1) : ((('h4000e7c8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomSymCalibOvlToClb                           = { [ (('h4000e7d0 - 'h4000d668) >> 1) : ((('h4000e7d0 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomAuxMeasResClbToOvl                         = { [ (('h4000e7d8 - 'h4000d668) >> 1) : ((('h4000e7d8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomCalibResClbToOvl                           = { [ (('h4000e7e0 - 'h4000d668) >> 1) : ((('h4000e7e0 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomSecDataKeysOtpToOvl                        = { [ (('h4000e7f8 - 'h4000d668) >> 1) : ((('h4000e7f8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomSecIdKeysOtpToOvl                          = { [ (('h4000e800 - 'h4000d668) >> 1) : ((('h4000e800 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomFmuOtpToOvl                                = { [ (('h4000e808 - 'h4000d668) >> 1) : ((('h4000e808 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomFmuOvlToClb                                = { [ (('h4000e810 - 'h4000d668) >> 1) : ((('h4000e810 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomFmuResHwsToOvl                             = { [ (('h4000e818 - 'h4000d668) >> 1) : ((('h4000e818 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomConfigFmuForLoDivSymVsSoc                  = { [ (('h4000e820 - 'h4000d668) >> 1) : ((('h4000e820 - 'h4000d668 + 'd32) >> 1) - 1) ] };
    bins SpuRomEnvdetMeasWithSoc                          = { [ (('h4000e840 - 'h4000d668) >> 1) : ((('h4000e840 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomCleOvlToHws                                = { [ (('h4000e858 - 'h4000d668) >> 1) : ((('h4000e858 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomCleHwsToOvl                                = { [ (('h4000e860 - 'h4000d668) >> 1) : ((('h4000e860 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomCleFllParams                               = { [ (('h4000e868 - 'h4000d668) >> 1) : ((('h4000e868 - 'h4000d668 + 'd28) >> 1) - 1) ] };
    bins SpuRomCopyCleAnalogctlForLcAuxIdacCalib          = { [ (('h4000e888 - 'h4000d668) >> 1) : ((('h4000e888 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomCopyCleAnalogctlForWkupThresholdCalib      = { [ (('h4000e890 - 'h4000d668) >> 1) : ((('h4000e890 - 'h4000d668 + 'd128) >> 1) - 1) ] };
    bins SpuRomCopyCleAnalogctlForLoVrefVbpCalib          = { [ (('h4000e910 - 'h4000d668) >> 1) : ((('h4000e910 - 'h4000d668 + 'd52) >> 1) - 1) ] };
    bins SpuRomCopyCleAnalogctlForDfCalib                 = { [ (('h4000e948 - 'h4000d668) >> 1) : ((('h4000e948 - 'h4000d668 + 'd16) >> 1) - 1) ] };
    bins SpuRomLoVrefVbpCalibRemoveSampling               = { [ (('h4000e958 - 'h4000d668) >> 1) : ((('h4000e958 - 'h4000d668 + 'd44) >> 1) - 1) ] };
    bins SpuRomSetVbpRxForCh39                            = { [ (('h4000e988 - 'h4000d668) >> 1) : ((('h4000e988 - 'h4000d668 + 'd36) >> 1) - 1) ] };
    bins SpuRomConfigFllForAuxMeas                        = { [ (('h4000e9b0 - 'h4000d668) >> 1) : ((('h4000e9b0 - 'h4000d668 + 'd32) >> 1) - 1) ] };
    bins SpuRomConfigFllForLoCalib                        = { [ (('h4000e9d0 - 'h4000d668) >> 1) : ((('h4000e9d0 - 'h4000d668 + 'd52) >> 1) - 1) ] };
    bins SpuRomConfigFllForSymCalib                       = { [ (('h4000ea08 - 'h4000d668) >> 1) : ((('h4000ea08 - 'h4000d668 + 'd32) >> 1) - 1) ] };
    bins SpuRomWaitFromOtp                                = { [ (('h4000ea28 - 'h4000d668) >> 1) : ((('h4000ea28 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomSetFlowManagerFsmCycleBeginInd0            = { [ (('h4000ea30 - 'h4000d668) >> 1) : ((('h4000ea30 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomSetFlowManagerFsmCycleBeginInd1            = { [ (('h4000ea38 - 'h4000d668) >> 1) : ((('h4000ea38 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomWkupStateCca                               = { [ (('h4000ea40 - 'h4000d668) >> 1) : ((('h4000ea40 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomWkupStateCh37                              = { [ (('h4000ea50 - 'h4000d668) >> 1) : ((('h4000ea50 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomWkupStateCh38                              = { [ (('h4000ea60 - 'h4000d668) >> 1) : ((('h4000ea60 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomWkupStateCh39                              = { [ (('h4000ea70 - 'h4000d668) >> 1) : ((('h4000ea70 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomSaveEaWkupTimers                           = { [ (('h4000ea80 - 'h4000d668) >> 1) : ((('h4000ea80 - 'h4000d668 + 'd40) >> 1) - 1) ] };
    bins SpuRomVddDig2VddAdbDisable                       = { [ (('h4000eaa8 - 'h4000d668) >> 1) : ((('h4000eaa8 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomVddDig2VddAdbEnable                        = { [ (('h4000eab0 - 'h4000d668) >> 1) : ((('h4000eab0 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomSetMaxEnvdetClkFreq                        = { [ (('h4000eab8 - 'h4000d668) >> 1) : ((('h4000eab8 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomSetMaxAttenuation                          = { [ (('h4000eac8 - 'h4000d668) >> 1) : ((('h4000eac8 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomSetMinAttenuation                          = { [ (('h4000ead8 - 'h4000d668) >> 1) : ((('h4000ead8 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomSetSlimLdoTrimForContWkup                  = { [ (('h4000eae0 - 'h4000d668) >> 1) : ((('h4000eae0 - 'h4000d668 + 'd40) >> 1) - 1) ] };
    bins SpuRomRestoreSlimLdoTrimAfterContWkup            = { [ (('h4000eb08 - 'h4000d668) >> 1) : ((('h4000eb08 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomSetPacketStructureInPacket                 = { [ (('h4000eb20 - 'h4000d668) >> 1) : ((('h4000eb20 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuCopyGroupID                                   = { [ (('h4000eb38 - 'h4000d668) >> 1) : ((('h4000eb38 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomInitializeUID                              = { [ (('h4000eb40 - 'h4000d668) >> 1) : ((('h4000eb40 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomCopyFlowVersionToPacketFromGnvm            = { [ (('h4000eb48 - 'h4000d668) >> 1) : ((('h4000eb48 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomUseMaxLcAuxFreq                            = { [ (('h4000eb58 - 'h4000d668) >> 1) : ((('h4000eb58 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomSetLcAuxFreqForTrng                        = { [ (('h4000eb60 - 'h4000d668) >> 1) : ((('h4000eb60 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomSetSymFreqForTrng                          = { [ (('h4000eb78 - 'h4000d668) >> 1) : ((('h4000eb78 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomCopyTrngToNonceSrr                         = { [ (('h4000eb90 - 'h4000d668) >> 1) : ((('h4000eb90 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomCopyTrngToAdvaSrr                          = { [ (('h4000eb98 - 'h4000d668) >> 1) : ((('h4000eb98 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomCopyTempEventCounterToGroupID              = { [ (('h4000eba0 - 'h4000d668) >> 1) : ((('h4000eba0 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomElevatorGearConfig                         = { [ (('h4000ebb8 - 'h4000d668) >> 1) : ((('h4000ebb8 - 'h4000d668 + 'd68) >> 1) - 1) ] };
    bins SpuRomDisableGearShiftTOExcptn                   = { [ (('h4000ec00 - 'h4000d668) >> 1) : ((('h4000ec00 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomHighGearConfig                             = { [ (('h4000ec18 - 'h4000d668) >> 1) : ((('h4000ec18 - 'h4000d668 + 'd108) >> 1) - 1) ] };
    bins SpuRomMidGearConfig                              = { [ (('h4000ec88 - 'h4000d668) >> 1) : ((('h4000ec88 - 'h4000d668 + 'd112) >> 1) - 1) ] };
    bins SpuRomPowerGearCheckGearReached                  = { [ (('h4000ecf8 - 'h4000d668) >> 1) : ((('h4000ecf8 - 'h4000d668 + 'd36) >> 1) - 1) ] };
    bins SpuRomPowerGearConfigHighGearSteadyState         = { [ (('h4000ed20 - 'h4000d668) >> 1) : ((('h4000ed20 - 'h4000d668 + 'd72) >> 1) - 1) ] };
    bins SpuRomPowerGearingExit                           = { [ (('h4000ed68 - 'h4000d668) >> 1) : ((('h4000ed68 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomPowerGearSetTimerForElevatorGear           = { [ (('h4000ed78 - 'h4000d668) >> 1) : ((('h4000ed78 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomPowerGearSetTimerForHighGear               = { [ (('h4000ed90 - 'h4000d668) >> 1) : ((('h4000ed90 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomPowerGearSetPowerGearingInd                = { [ (('h4000eda8 - 'h4000d668) >> 1) : ((('h4000eda8 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomPowerGearClearPowerGearingInd              = { [ (('h4000edb0 - 'h4000d668) >> 1) : ((('h4000edb0 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomPowerGearSetFastHarvester                  = { [ (('h4000edb8 - 'h4000d668) >> 1) : ((('h4000edb8 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomPowerGearSetSlowHarvester                  = { [ (('h4000edc8 - 'h4000d668) >> 1) : ((('h4000edc8 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins setFmuInitMask                                   = { [ (('h4000edd8 - 'h4000d668) >> 1) : ((('h4000edd8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomFixControl                                 = { [ (('h4000ede0 - 'h4000d668) >> 1) : ((('h4000ede0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomFixTimer                                   = { [ (('h4000edf8 - 'h4000d668) >> 1) : ((('h4000edf8 - 'h4000d668 + 'd16) >> 1) - 1) ] };
    bins spuRomEvent0FixControl                           = { [ (('h4000ee08 - 'h4000d668) >> 1) : ((('h4000ee08 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent0FixTimer                             = { [ (('h4000ee10 - 'h4000d668) >> 1) : ((('h4000ee10 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent1FixControl                           = { [ (('h4000ee18 - 'h4000d668) >> 1) : ((('h4000ee18 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent1FixTimer                             = { [ (('h4000ee20 - 'h4000d668) >> 1) : ((('h4000ee20 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent2FixControl                           = { [ (('h4000ee28 - 'h4000d668) >> 1) : ((('h4000ee28 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent2FixTimer                             = { [ (('h4000ee30 - 'h4000d668) >> 1) : ((('h4000ee30 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent3FixControl                           = { [ (('h4000ee38 - 'h4000d668) >> 1) : ((('h4000ee38 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent3FixTimer                             = { [ (('h4000ee40 - 'h4000d668) >> 1) : ((('h4000ee40 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent4FixControl                           = { [ (('h4000ee48 - 'h4000d668) >> 1) : ((('h4000ee48 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent4FixTimer                             = { [ (('h4000ee50 - 'h4000d668) >> 1) : ((('h4000ee50 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent5FixControl                           = { [ (('h4000ee58 - 'h4000d668) >> 1) : ((('h4000ee58 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent5FixTimer                             = { [ (('h4000ee60 - 'h4000d668) >> 1) : ((('h4000ee60 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent6FixControl                           = { [ (('h4000ee68 - 'h4000d668) >> 1) : ((('h4000ee68 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent6FixTimer                             = { [ (('h4000ee70 - 'h4000d668) >> 1) : ((('h4000ee70 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent7FixControl                           = { [ (('h4000ee78 - 'h4000d668) >> 1) : ((('h4000ee78 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent7FixTimer                             = { [ (('h4000ee80 - 'h4000d668) >> 1) : ((('h4000ee80 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent8FixControl                           = { [ (('h4000ee88 - 'h4000d668) >> 1) : ((('h4000ee88 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent8FixTimer                             = { [ (('h4000ee90 - 'h4000d668) >> 1) : ((('h4000ee90 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent9FixControl                           = { [ (('h4000ee98 - 'h4000d668) >> 1) : ((('h4000ee98 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent9FixTimer                             = { [ (('h4000eea0 - 'h4000d668) >> 1) : ((('h4000eea0 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent10FixControl                          = { [ (('h4000eea8 - 'h4000d668) >> 1) : ((('h4000eea8 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent10FixTimer                            = { [ (('h4000eeb0 - 'h4000d668) >> 1) : ((('h4000eeb0 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent11FixControl                          = { [ (('h4000eeb8 - 'h4000d668) >> 1) : ((('h4000eeb8 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent11FixTimer                            = { [ (('h4000eec0 - 'h4000d668) >> 1) : ((('h4000eec0 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent12FixControl                          = { [ (('h4000eec8 - 'h4000d668) >> 1) : ((('h4000eec8 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent12FixTimer                            = { [ (('h4000eed0 - 'h4000d668) >> 1) : ((('h4000eed0 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent13FixControl                          = { [ (('h4000eed8 - 'h4000d668) >> 1) : ((('h4000eed8 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent13FixTimer                            = { [ (('h4000eee0 - 'h4000d668) >> 1) : ((('h4000eee0 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent14FixControl                          = { [ (('h4000eee8 - 'h4000d668) >> 1) : ((('h4000eee8 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent14FixTimer                            = { [ (('h4000eef0 - 'h4000d668) >> 1) : ((('h4000eef0 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent15FixControl                          = { [ (('h4000eef8 - 'h4000d668) >> 1) : ((('h4000eef8 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomEvent15FixTimer                            = { [ (('h4000ef00 - 'h4000d668) >> 1) : ((('h4000ef00 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins spuRomTurnOffMss                                 = { [ (('h4000ef08 - 'h4000d668) >> 1) : ((('h4000ef08 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins spuRomTurnOffRadio                               = { [ (('h4000ef18 - 'h4000d668) >> 1) : ((('h4000ef18 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomRtcSocMeas                                 = { [ (('h4000ef30 - 'h4000d668) >> 1) : ((('h4000ef30 - 'h4000d668 + 'd52) >> 1) - 1) ] };
    bins SpuRomVstartCalibInit                            = { [ (('h4000ef68 - 'h4000d668) >> 1) : ((('h4000ef68 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomTestSecSetup                               = { [ (('h4000ef80 - 'h4000d668) >> 1) : ((('h4000ef80 - 'h4000d668 + 'd60) >> 1) - 1) ] };
    bins SpuRomByteAccessSRR                              = { [ (('h4000efc0 - 'h4000d668) >> 1) : ((('h4000efc0 - 'h4000d668 + 'd28) >> 1) - 1) ] };
    bins SpuRomPopulateRadioHws                           = { [ (('h4000efe0 - 'h4000d668) >> 1) : ((('h4000efe0 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomSymMeasLcRadioInit                         = { [ (('h4000efe8 - 'h4000d668) >> 1) : ((('h4000efe8 - 'h4000d668 + 'd80) >> 1) - 1) ] };
    bins SpuRomRadioModeSymMeasLc                         = { [ (('h4000f038 - 'h4000d668) >> 1) : ((('h4000f038 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomLcauxIdacCalibInit                         = { [ (('h4000f048 - 'h4000d668) >> 1) : ((('h4000f048 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomUnSetFirstCycleCalibIter                   = { [ (('h4000f060 - 'h4000d668) >> 1) : ((('h4000f060 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomBasicFlowCopyClbCfgOTPToIsp                = { [ (('h4000f068 - 'h4000d668) >> 1) : ((('h4000f068 - 'h4000d668 + 'd36) >> 1) - 1) ] };
    bins SpuRomBasicFlowAuxMeasCfgIspToOvl                = { [ (('h4000f090 - 'h4000d668) >> 1) : ((('h4000f090 - 'h4000d668 + 'd16) >> 1) - 1) ] };
    bins SpuRomBasicFlowLoClbIspToOvl                     = { [ (('h4000f0a0 - 'h4000d668) >> 1) : ((('h4000f0a0 - 'h4000d668 + 'd24) >> 1) - 1) ] };
    bins SpuRomBasicFlowSymClbIspToOvl                    = { [ (('h4000f0b8 - 'h4000d668) >> 1) : ((('h4000f0b8 - 'h4000d668 + 'd16) >> 1) - 1) ] };
    bins SpuRomBasicFlowPreparePacketWithConst            = { [ (('h4000f0c8 - 'h4000d668) >> 1) : ((('h4000f0c8 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomBasicFlowPreparePacketWithSec              = { [ (('h4000f0e0 - 'h4000d668) >> 1) : ((('h4000f0e0 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomBasicFlowKeepOtpShutOffEn                  = { [ (('h4000f0e8 - 'h4000d668) >> 1) : ((('h4000f0e8 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomBasicFlowSpuNOP                            = { [ (('h4000f0f0 - 'h4000d668) >> 1) : ((('h4000f0f0 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins RET_init_from_GNVM                               = { [ (('h4000f0f8 - 'h4000d668) >> 1) : ((('h4000f0f8 - 'h4000d668 + 'd64) >> 1) - 1) ] };
    bins CLB_init_from_GNVM                               = { [ (('h4000f138 - 'h4000d668) >> 1) : ((('h4000f138 - 'h4000d668 + 'd28) >> 1) - 1) ] };
    bins SpuRomFirstBootInit                              = { [ (('h4000f158 - 'h4000d668) >> 1) : ((('h4000f158 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins spuRomInitFromGnvm                               = { [ (('h4000f168 - 'h4000d668) >> 1) : ((('h4000f168 - 'h4000d668 + 'd64) >> 1) - 1) ] };
    bins SpuRomSetWuParamsForTestModeWU                   = { [ (('h4000f1a8 - 'h4000d668) >> 1) : ((('h4000f1a8 - 'h4000d668 + 'd64) >> 1) - 1) ] };
    bins SpuRomSetAueMeasTimeTo2                          = { [ (('h4000f1e8 - 'h4000d668) >> 1) : ((('h4000f1e8 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomTestModeSetWuState12                       = { [ (('h4000f1f8 - 'h4000d668) >> 1) : ((('h4000f1f8 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomTestModeSetWuState14                       = { [ (('h4000f208 - 'h4000d668) >> 1) : ((('h4000f208 - 'h4000d668 + 'd12) >> 1) - 1) ] };
    bins SpuRomForceReset                                 = { [ (('h4000f218 - 'h4000d668) >> 1) : ((('h4000f218 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomDisableSoftAWDT                            = { [ (('h4000f220 - 'h4000d668) >> 1) : ((('h4000f220 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomHwsRegistersInitFromGnvm                   = { [ (('h4000f228 - 'h4000d668) >> 1) : ((('h4000f228 - 'h4000d668 + 'd20) >> 1) - 1) ] };
    bins SpuRomHwsHrrInitFromGnvm                         = { [ (('h4000f240 - 'h4000d668) >> 1) : ((('h4000f240 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomIspSrrInitFromGnvm                         = { [ (('h4000f248 - 'h4000d668) >> 1) : ((('h4000f248 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuRomAuxMeasAndCalibOverlayInitFromGnvm         = { [ (('h4000f250 - 'h4000d668) >> 1) : ((('h4000f250 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomSecAndTxOverlayInitFromGnvm                = { [ (('h4000f258 - 'h4000d668) >> 1) : ((('h4000f258 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomFlowManagerAndPowerupOverlayInitFromGnvm   = { [ (('h4000f260 - 'h4000d668) >> 1) : ((('h4000f260 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomPowerGearingOverlayInitFromGnvm            = { [ (('h4000f268 - 'h4000d668) >> 1) : ((('h4000f268 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomLcAuxIdacCalibOverlayInitFromGnvm          = { [ (('h4000f270 - 'h4000d668) >> 1) : ((('h4000f270 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomWkupThresholdCalibOverlayInitFromGnvm      = { [ (('h4000f278 - 'h4000d668) >> 1) : ((('h4000f278 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomLoVrefVbpCalibOverlayInitFromGnvm          = { [ (('h4000f280 - 'h4000d668) >> 1) : ((('h4000f280 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomDfCalibOverlayInitFromGnvm                 = { [ (('h4000f288 - 'h4000d668) >> 1) : ((('h4000f288 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomSensingOverlayInitFromGnvm                 = { [ (('h4000f290 - 'h4000d668) >> 1) : ((('h4000f290 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomTempPolyCoeffOverlayInitFromGnvm           = { [ (('h4000f298 - 'h4000d668) >> 1) : ((('h4000f298 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomAuxMeasVsTempCoeffOverlayInitFromGnvm      = { [ (('h4000f2a0 - 'h4000d668) >> 1) : ((('h4000f2a0 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomTestModeOverlayInitFromGnvm                = { [ (('h4000f2a8 - 'h4000d668) >> 1) : ((('h4000f2a8 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomSystemClksMeasOverlayInitFromGnvm          = { [ (('h4000f2b0 - 'h4000d668) >> 1) : ((('h4000f2b0 - 'h4000d668 + 'd4) >> 1) - 1) ] };
    bins SpuRomClbRegistersInitFromGnvm                   = { [ (('h4000f2b8 - 'h4000d668) >> 1) : ((('h4000f2b8 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuNvmTestFunction                               = { [ (('h40010c00 - 'h4000d668) >> 1) : ((('h40010c00 - 'h4000d668 + 'd8) >> 1) - 1) ] };
    bins SpuNvmTestFunction2                              = { [ (('h40010c08 - 'h4000d668) >> 1) : ((('h40010c08 - 'h4000d668 + 'd12) >> 1) - 1) ] };