    bins _start                                                       = { [ (('h40000000 - 'h40000000) >> 1) : ((('h40000000 - 'h40000000 + 'd36) >> 1) - 1) ] };
    bins rom_index                                                    = { [ (('h40000030 - 'h40000000) >> 1) : ((('h40000030 - 'h40000000 + 'd4) >> 1) - 1) ] };
    bins FlowExceptionHandler                                         = { [ (('h40000040 - 'h40000000) >> 1) : ((('h40000040 - 'h40000000 + 'd36) >> 1) - 1) ] };
    bins MachineTrapEntry                                             = { [ (('h40000080 - 'h40000000) >> 1) : ((('h40000080 - 'h40000000 + 'd26) >> 1) - 1) ] };
    bins McuRomDma                                                    = { [ (('h40000210 - 'h40000000) >> 1) : ((('h40000210 - 'h40000000 + 'd50) >> 1) - 1) ] };
    bins McuRomOtpProgDma                                             = { [ (('h40000248 - 'h40000000) >> 1) : ((('h40000248 - 'h40000000 + 'd112) >> 1) - 1) ] };
    bins McuRomOtpCompare                                             = { [ (('h400002b8 - 'h40000000) >> 1) : ((('h400002b8 - 'h40000000 + 'd40) >> 1) - 1) ] };
    bins McuRomSimpleDma                                              = { [ (('h400002e0 - 'h40000000) >> 1) : ((('h400002e0 - 'h40000000 + 'd54) >> 1) - 1) ] };
    bins McuRomVerifyDma                                              = { [ (('h40000318 - 'h40000000) >> 1) : ((('h40000318 - 'h40000000 + 'd90) >> 1) - 1) ] };
    bins McuRomVerifyCrc                                              = { [ (('h40000378 - 'h40000000) >> 1) : ((('h40000378 - 'h40000000 + 'd42) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForTxLv                         = { [ (('h400003a8 - 'h40000000) >> 1) : ((('h400003a8 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForTxLv                         = { [ (('h400003e8 - 'h40000000) >> 1) : ((('h400003e8 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForLoCalibLv                    = { [ (('h400003f8 - 'h40000000) >> 1) : ((('h400003f8 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForLoCalibLv                    = { [ (('h40000438 - 'h40000000) >> 1) : ((('h40000438 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForMeasureLv                    = { [ (('h40000448 - 'h40000000) >> 1) : ((('h40000448 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForMeasureLv                    = { [ (('h40000488 - 'h40000000) >> 1) : ((('h40000488 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForSymCalibLv                   = { [ (('h40000498 - 'h40000000) >> 1) : ((('h40000498 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForSymCalibLv                   = { [ (('h400004d8 - 'h40000000) >> 1) : ((('h400004d8 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForTxHv                         = { [ (('h400004e8 - 'h40000000) >> 1) : ((('h400004e8 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForTxHv                         = { [ (('h40000528 - 'h40000000) >> 1) : ((('h40000528 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForLoCalibHv                    = { [ (('h40000538 - 'h40000000) >> 1) : ((('h40000538 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForLoCalibHv                    = { [ (('h40000578 - 'h40000000) >> 1) : ((('h40000578 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForMeasureHv                    = { [ (('h40000588 - 'h40000000) >> 1) : ((('h40000588 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForMeasureHv                    = { [ (('h400005c8 - 'h40000000) >> 1) : ((('h400005c8 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForSymCalibHv                   = { [ (('h400005d8 - 'h40000000) >> 1) : ((('h400005d8 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForSymCalibHv                   = { [ (('h40000618 - 'h40000000) >> 1) : ((('h40000618 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForTempsensLv                   = { [ (('h40000628 - 'h40000000) >> 1) : ((('h40000628 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForTempsensLv                   = { [ (('h40000668 - 'h40000000) >> 1) : ((('h40000668 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForMeasureLC                    = { [ (('h40000678 - 'h40000000) >> 1) : ((('h40000678 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForMeasureLC                    = { [ (('h400006b8 - 'h40000000) >> 1) : ((('h400006b8 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForrcSensCap                    = { [ (('h400006c8 - 'h40000000) >> 1) : ((('h400006c8 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForrcSensCap                    = { [ (('h40000708 - 'h40000000) >> 1) : ((('h40000708 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForrcSensRes                    = { [ (('h40000718 - 'h40000000) >> 1) : ((('h40000718 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForrcSensRes                    = { [ (('h40000758 - 'h40000000) >> 1) : ((('h40000758 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForLoDivSymLv                   = { [ (('h40000768 - 'h40000000) >> 1) : ((('h40000768 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetModeTableAddressForLoDivSymHv                   = { [ (('h40000778 - 'h40000000) >> 1) : ((('h40000778 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForLoDivSymLv                   = { [ (('h40000788 - 'h40000000) >> 1) : ((('h40000788 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins mcuRomFlowSetInitTableAddressForLoDivSymHv                   = { [ (('h400007c8 - 'h40000000) >> 1) : ((('h400007c8 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins RomSetBatteryAndHpmModes                                     = { [ (('h40000808 - 'h40000000) >> 1) : ((('h40000808 - 'h40000000 + 'd88) >> 1) - 1) ] };
    bins CalibAndTxFsmSetTxoRxoPerPowerMode                           = { [ (('h40000860 - 'h40000000) >> 1) : ((('h40000860 - 'h40000000 + 'd94) >> 1) - 1) ] };
    bins CalcTempRange                                                = { [ (('h400008c0 - 'h40000000) >> 1) : ((('h400008c0 - 'h40000000 + 'd144) >> 1) - 1) ] };
    bins TempCompAnalogControl                                        = { [ (('h40000950 - 'h40000000) >> 1) : ((('h40000950 - 'h40000000 + 'd110) >> 1) - 1) ] };
    bins TempCompAnalogControlWithoutUpdatingTempCompVector           = { [ (('h400009c0 - 'h40000000) >> 1) : ((('h400009c0 - 'h40000000 + 'd90) >> 1) - 1) ] };
    bins TempCompAnalogRguWsContext0ParamsSetOffsets                  = { [ (('h40000a20 - 'h40000000) >> 1) : ((('h40000a20 - 'h40000000 + 'd90) >> 1) - 1) ] };
    bins TempCompAnalogRguWsContext1ParamsSetOffsets                  = { [ (('h40000a80 - 'h40000000) >> 1) : ((('h40000a80 - 'h40000000 + 'd90) >> 1) - 1) ] };
    bins TempCompAnalogRguDynClbAndTempLoopContextParamsSetOffsets    = { [ (('h40000ae0 - 'h40000000) >> 1) : ((('h40000ae0 - 'h40000000 + 'd146) >> 1) - 1) ] };
    bins TempCompAnalogHrrAndDrrShadowParamsSetOffsets                = { [ (('h40000b78 - 'h40000000) >> 1) : ((('h40000b78 - 'h40000000 + 'd146) >> 1) - 1) ] };
    bins TempCompAnalogRguWsContext0ParamsExecute                     = { [ (('h40000c10 - 'h40000000) >> 1) : ((('h40000c10 - 'h40000000 + 'd402) >> 1) - 1) ] };
    bins TempCompAnalogRguWsContext1ParamsExecute                     = { [ (('h40000da8 - 'h40000000) >> 1) : ((('h40000da8 - 'h40000000 + 'd466) >> 1) - 1) ] };
    bins TempCompAnalogRguDynClbAndTempLoopContextParamsExecute       = { [ (('h40000f80 - 'h40000000) >> 1) : ((('h40000f80 - 'h40000000 + 'd526) >> 1) - 1) ] };
    bins TempCompSlimLdo                                              = { [ (('h40001190 - 'h40000000) >> 1) : ((('h40001190 - 'h40000000 + 'd206) >> 1) - 1) ] };
    bins TempCompAnalogHrrAndDrrShadowParamsExecute                   = { [ (('h40001260 - 'h40000000) >> 1) : ((('h40001260 - 'h40000000 + 'd550) >> 1) - 1) ] };
    bins TempCompEnvdetClkCoarse                                      = { [ (('h40001488 - 'h40000000) >> 1) : ((('h40001488 - 'h40000000 + 'd106) >> 1) - 1) ] };
    bins TempCompDigLdo                                               = { [ (('h400014f8 - 'h40000000) >> 1) : ((('h400014f8 - 'h40000000 + 'd96) >> 1) - 1) ] };
    bins TempCompActiveClkTrim                                        = { [ (('h40001558 - 'h40000000) >> 1) : ((('h40001558 - 'h40000000 + 'd96) >> 1) - 1) ] };
    bins TempCompRtcClkTrim                                           = { [ (('h400015b8 - 'h40000000) >> 1) : ((('h400015b8 - 'h40000000 + 'd106) >> 1) - 1) ] };
    bins CalcAuxFreqCompFactor                                        = { [ (('h40001628 - 'h40000000) >> 1) : ((('h40001628 - 'h40000000 + 'd24) >> 1) - 1) ] };
    bins EstAuxFreqForTemperatureAndHypothesis                        = { [ (('h40001640 - 'h40000000) >> 1) : ((('h40001640 - 'h40000000 + 'd298) >> 1) - 1) ] };
    bins McuRomResetCleOvl                                            = { [ (('h40001770 - 'h40000000) >> 1) : ((('h40001770 - 'h40000000 + 'd14) >> 1) - 1) ] };
    bins CtlCalibInit                                                 = { [ (('h40001780 - 'h40000000) >> 1) : ((('h40001780 - 'h40000000 + 'd78) >> 1) - 1) ] };
    bins CtlCalibResetCoarseStepSize                                  = { [ (('h400017d0 - 'h40000000) >> 1) : ((('h400017d0 - 'h40000000 + 'd20) >> 1) - 1) ] };
    bins CtlCalibUpdateControls                                       = { [ (('h400017e8 - 'h40000000) >> 1) : ((('h400017e8 - 'h40000000 + 'd104) >> 1) - 1) ] };
    bins CtlCalibFsm                                                  = { [ (('h40001850 - 'h40000000) >> 1) : ((('h40001850 - 'h40000000 + 'd398) >> 1) - 1) ] };
    bins CtlCalibIncStateUponSignalToggle                             = { [ (('h400019e0 - 'h40000000) >> 1) : ((('h400019e0 - 'h40000000 + 'd44) >> 1) - 1) ] };
    bins CleCheckIfMaxStepReached                                     = { [ (('h40001a10 - 'h40000000) >> 1) : ((('h40001a10 - 'h40000000 + 'd66) >> 1) - 1) ] };
    bins LoVrefVbpCalibSaveCurrConfigForDebugData                     = { [ (('h40001a58 - 'h40000000) >> 1) : ((('h40001a58 - 'h40000000 + 'd106) >> 1) - 1) ] };
    bins LoVrefVbpCalibCleInit                                        = { [ (('h40001ac8 - 'h40000000) >> 1) : ((('h40001ac8 - 'h40000000 + 'd242) >> 1) - 1) ] };
    bins LoVrefVbpCalibCleOverflow                                    = { [ (('h40001bc0 - 'h40000000) >> 1) : ((('h40001bc0 - 'h40000000 + 'd218) >> 1) - 1) ] };
    bins LoVrefVbpCalibSetCoarseStepSize                              = { [ (('h40001ca0 - 'h40000000) >> 1) : ((('h40001ca0 - 'h40000000 + 'd94) >> 1) - 1) ] };
    bins LoVrefVbpCalibSetVrefTxField                                 = { [ (('h40001d00 - 'h40000000) >> 1) : ((('h40001d00 - 'h40000000 + 'd34) >> 1) - 1) ] };
    bins LoVrefVbpCalibSetVrefRxField                                 = { [ (('h40001d28 - 'h40000000) >> 1) : ((('h40001d28 - 'h40000000 + 'd34) >> 1) - 1) ] };
    bins LoVrefVbpCalibGetVrefTxField                                 = { [ (('h40001d50 - 'h40000000) >> 1) : ((('h40001d50 - 'h40000000 + 'd42) >> 1) - 1) ] };
    bins LoVrefVbpCalibGetVrefRxField                                 = { [ (('h40001d80 - 'h40000000) >> 1) : ((('h40001d80 - 'h40000000 + 'd42) >> 1) - 1) ] };
    bins LoVrefVbpCalibEnsureOscillationUponDone                      = { [ (('h40001db0 - 'h40000000) >> 1) : ((('h40001db0 - 'h40000000 + 'd70) >> 1) - 1) ] };
    bins LoVrefVbpCalibSaveControls                                   = { [ (('h40001df8 - 'h40000000) >> 1) : ((('h40001df8 - 'h40000000 + 'd206) >> 1) - 1) ] };
    bins LoVrefVbpCalibRestoreControls                                = { [ (('h40001ec8 - 'h40000000) >> 1) : ((('h40001ec8 - 'h40000000 + 'd198) >> 1) - 1) ] };
    bins LoVrefVbpCalibFinalizeTxControls                             = { [ (('h40001f90 - 'h40000000) >> 1) : ((('h40001f90 - 'h40000000 + 'd178) >> 1) - 1) ] };
    bins LoVrefVbpCalibFinalizeRxControls                             = { [ (('h40002048 - 'h40000000) >> 1) : ((('h40002048 - 'h40000000 + 'd176) >> 1) - 1) ] };
    bins LoVrefVbpCalibFinalizeControls                               = { [ (('h400020f8 - 'h40000000) >> 1) : ((('h400020f8 - 'h40000000 + 'd44) >> 1) - 1) ] };
    bins LoVrefVbpCalibResetControlsToGnvm                            = { [ (('h40002128 - 'h40000000) >> 1) : ((('h40002128 - 'h40000000 + 'd250) >> 1) - 1) ] };
    bins LoVrefVbpCalibCopyTxCtrlsToRxCtrls                           = { [ (('h40002228 - 'h40000000) >> 1) : ((('h40002228 - 'h40000000 + 'd78) >> 1) - 1) ] };
    bins LoVrefVbpCalibUpdateControlsForVerifUponConsecBadCalibs      = { [ (('h40002278 - 'h40000000) >> 1) : ((('h40002278 - 'h40000000 + 'd84) >> 1) - 1) ] };
    bins LoVrefVbpCalibUpdateBadCalibCtr                              = { [ (('h400022d0 - 'h40000000) >> 1) : ((('h400022d0 - 'h40000000 + 'd74) >> 1) - 1) ] };
    bins LoVrefVbpCalibCheckConsecutiveBeacons                        = { [ (('h40002320 - 'h40000000) >> 1) : ((('h40002320 - 'h40000000 + 'd158) >> 1) - 1) ] };
    bins LoVrefVbpCalibUseLcAuxForVerification                        = { [ (('h400023c0 - 'h40000000) >> 1) : ((('h400023c0 - 'h40000000 + 'd52) >> 1) - 1) ] };
    bins LcAuxCalibEnsureOscillationUponDone                          = { [ (('h400023f8 - 'h40000000) >> 1) : ((('h400023f8 - 'h40000000 + 'd74) >> 1) - 1) ] };
    bins LcAuxCalibResetControlsToGnvm                                = { [ (('h40002448 - 'h40000000) >> 1) : ((('h40002448 - 'h40000000 + 'd22) >> 1) - 1) ] };
    bins LcAuxCalibSaveCurrConfigForDebugData                         = { [ (('h40002460 - 'h40000000) >> 1) : ((('h40002460 - 'h40000000 + 'd42) >> 1) - 1) ] };
    bins DfCalibSaveCurrConfigForDebugData                            = { [ (('h40002490 - 'h40000000) >> 1) : ((('h40002490 - 'h40000000 + 'd42) >> 1) - 1) ] };
    bins DfCalibCleCalcSprinklerEfineStep                             = { [ (('h400024c0 - 'h40000000) >> 1) : ((('h400024c0 - 'h40000000 + 'd50) >> 1) - 1) ] };
    bins PrepareFirstDfMeas                                           = { [ (('h400024f8 - 'h40000000) >> 1) : ((('h400024f8 - 'h40000000 + 'd194) >> 1) - 1) ] };
    bins RomSetTxDfAndSprinklerForSmallStepEfine                      = { [ (('h400025c0 - 'h40000000) >> 1) : ((('h400025c0 - 'h40000000 + 'd62) >> 1) - 1) ] };
    bins RomSetTxDfAndSprinklerForNormalStepEfine                     = { [ (('h40002600 - 'h40000000) >> 1) : ((('h40002600 - 'h40000000 + 'd62) >> 1) - 1) ] };
    bins BleFreqMhzToChIdx                                            = { [ (('h40002640 - 'h40000000) >> 1) : ((('h40002640 - 'h40000000 + 'd78) >> 1) - 1) ] };
    bins BleChIdxToFreqMhz                                            = { [ (('h40002690 - 'h40000000) >> 1) : ((('h40002690 - 'h40000000 + 'd84) >> 1) - 1) ] };
    bins CalcCwScalerFromGivenBleChIdx                                = { [ (('h400026e8 - 'h40000000) >> 1) : ((('h400026e8 - 'h40000000 + 'd118) >> 1) - 1) ] };
    bins CalcLoDivSymDivRatioFromGivenBleChIdx                        = { [ (('h40002760 - 'h40000000) >> 1) : ((('h40002760 - 'h40000000 + 'd152) >> 1) - 1) ] };
    bins McuRomAuxMeasPrepare                                         = { [ (('h400027f8 - 'h40000000) >> 1) : ((('h400027f8 - 'h40000000 + 'd666) >> 1) - 1) ] };
    bins McuRomRxSweepPreProcessing                                   = { [ (('h40002a98 - 'h40000000) >> 1) : ((('h40002a98 - 'h40000000 + 'd324) >> 1) - 1) ] };
    bins McuRomRxSweepPostProcessing                                  = { [ (('h40002be0 - 'h40000000) >> 1) : ((('h40002be0 - 'h40000000 + 'd316) >> 1) - 1) ] };
    bins CalibAndTxFsmAuxMeas                                         = { [ (('h40002d20 - 'h40000000) >> 1) : ((('h40002d20 - 'h40000000 + 'd4) >> 1) - 1) ] };
    bins CalibAndTxFsmUpdateNrgdetDurationThr                         = { [ (('h40002d28 - 'h40000000) >> 1) : ((('h40002d28 - 'h40000000 + 'd152) >> 1) - 1) ] };
    bins CalibAndTxFsmCheckGoodAuxMeas                                = { [ (('h40002dc0 - 'h40000000) >> 1) : ((('h40002dc0 - 'h40000000 + 'd492) >> 1) - 1) ] };
    bins CalibAndTxFsmNoGoodAuxMeas                                   = { [ (('h40002fb0 - 'h40000000) >> 1) : ((('h40002fb0 - 'h40000000 + 'd178) >> 1) - 1) ] };
    bins CalibAndTxCheckDiscardRxSweep                                = { [ (('h40003068 - 'h40000000) >> 1) : ((('h40003068 - 'h40000000 + 'd162) >> 1) - 1) ] };
    bins McuRomAuxMeasPostProcessing                                  = { [ (('h40003110 - 'h40000000) >> 1) : ((('h40003110 - 'h40000000 + 'd294) >> 1) - 1) ] };
    bins CalibAndTxFsmLoTxRxCalib                                     = { [ (('h40003238 - 'h40000000) >> 1) : ((('h40003238 - 'h40000000 + 'd108) >> 1) - 1) ] };
    bins RomSetSprinklerDCO                                           = { [ (('h400032a8 - 'h40000000) >> 1) : ((('h400032a8 - 'h40000000 + 'd264) >> 1) - 1) ] };
    bins McuRomSetMaxTimeSprinkler                                    = { [ (('h400033b0 - 'h40000000) >> 1) : ((('h400033b0 - 'h40000000 + 'd154) >> 1) - 1) ] };
    bins McuRomSetMaxFreqSprinkler                                    = { [ (('h40003450 - 'h40000000) >> 1) : ((('h40003450 - 'h40000000 + 'd108) >> 1) - 1) ] };
    bins McuRomSetChannelSprinkler                                    = { [ (('h400034c0 - 'h40000000) >> 1) : ((('h400034c0 - 'h40000000 + 'd204) >> 1) - 1) ] };
    bins McuRomRestoreParamsUponTxSprinklerDone                       = { [ (('h40003590 - 'h40000000) >> 1) : ((('h40003590 - 'h40000000 + 'd234) >> 1) - 1) ] };
    bins McuRomMiniRxChooseHarvesterFlow                              = { [ (('h40003680 - 'h40000000) >> 1) : ((('h40003680 - 'h40000000 + 'd162) >> 1) - 1) ] };
    bins McuRomMiniRxChooseBle5FreqConfig                             = { [ (('h40003728 - 'h40000000) >> 1) : ((('h40003728 - 'h40000000 + 'd88) >> 1) - 1) ] };
    bins McuRomMiniRxChooseBle5PacketsConfig                          = { [ (('h40003780 - 'h40000000) >> 1) : ((('h40003780 - 'h40000000 + 'd66) >> 1) - 1) ] };
    bins McuRomMiniRxChooseHarvesterTypeConfig                        = { [ (('h400037c8 - 'h40000000) >> 1) : ((('h400037c8 - 'h40000000 + 'd34) >> 1) - 1) ] };
    bins McuRomMiniRxChooseBle5SymbolRateConfig                       = { [ (('h400037f0 - 'h40000000) >> 1) : ((('h400037f0 - 'h40000000 + 'd36) >> 1) - 1) ] };
    bins McuRomMiniRxChooseGearAndLoPmConfig                          = { [ (('h40003818 - 'h40000000) >> 1) : ((('h40003818 - 'h40000000 + 'd44) >> 1) - 1) ] };
    bins McuRomMiniRxForceVrefVbpConfig                               = { [ (('h40003848 - 'h40000000) >> 1) : ((('h40003848 - 'h40000000 + 'd438) >> 1) - 1) ] };
    bins McuRomMiniRxScanLoDcoConfig                                  = { [ (('h40003a00 - 'h40000000) >> 1) : ((('h40003a00 - 'h40000000 + 'd184) >> 1) - 1) ] };
    bins McuRomMiniRxSub1gHarvSwitchConfig                            = { [ (('h40003ab8 - 'h40000000) >> 1) : ((('h40003ab8 - 'h40000000 + 'd14) >> 1) - 1) ] };
    bins FmuFilter                                                    = { [ (('h40003ac8 - 'h40000000) >> 1) : ((('h40003ac8 - 'h40000000 + 'd70) >> 1) - 1) ] };
    bins FmuSetNumCycles                                              = { [ (('h40003b10 - 'h40000000) >> 1) : ((('h40003b10 - 'h40000000 + 'd26) >> 1) - 1) ] };
    bins MeasureClockFreqHz                                           = { [ (('h40003b30 - 'h40000000) >> 1) : ((('h40003b30 - 'h40000000 + 'd88) >> 1) - 1) ] };
    bins WkupCalibInit                                                = { [ (('h40003b88 - 'h40000000) >> 1) : ((('h40003b88 - 'h40000000 + 'd72) >> 1) - 1) ] };
    bins WkupCalibRestoreConfigUponCalibDone                          = { [ (('h40003bd0 - 'h40000000) >> 1) : ((('h40003bd0 - 'h40000000 + 'd142) >> 1) - 1) ] };
    bins WkupLowSensitivityCalibSetThreshold                          = { [ (('h40003c60 - 'h40000000) >> 1) : ((('h40003c60 - 'h40000000 + 'd100) >> 1) - 1) ] };
    bins WkupHighSensitivityCalibSetThreshold                         = { [ (('h40003cc8 - 'h40000000) >> 1) : ((('h40003cc8 - 'h40000000 + 'd156) >> 1) - 1) ] };
    bins WkupSample                                                   = { [ (('h40003d68 - 'h40000000) >> 1) : ((('h40003d68 - 'h40000000 + 'd246) >> 1) - 1) ] };
    bins RomSetWkupSensitivity                                        = { [ (('h40003e60 - 'h40000000) >> 1) : ((('h40003e60 - 'h40000000 + 'd100) >> 1) - 1) ] };
    bins WkupCalibCleInit                                             = { [ (('h40003ec8 - 'h40000000) >> 1) : ((('h40003ec8 - 'h40000000 + 'd250) >> 1) - 1) ] };
    bins WkupCalibSaveControls                                        = { [ (('h40003fc8 - 'h40000000) >> 1) : ((('h40003fc8 - 'h40000000 + 'd142) >> 1) - 1) ] };
    bins WkupCalibRestoreControls                                     = { [ (('h40004058 - 'h40000000) >> 1) : ((('h40004058 - 'h40000000 + 'd86) >> 1) - 1) ] };
    bins WkupCalibCleOverflow                                         = { [ (('h400040b0 - 'h40000000) >> 1) : ((('h400040b0 - 'h40000000 + 'd200) >> 1) - 1) ] };
    bins WkupCalibSaveCurrConfigForDebugData                          = { [ (('h40004178 - 'h40000000) >> 1) : ((('h40004178 - 'h40000000 + 'd130) >> 1) - 1) ] };
    bins WkupLowSensitivityCalibInit                                  = { [ (('h40004200 - 'h40000000) >> 1) : ((('h40004200 - 'h40000000 + 'd118) >> 1) - 1) ] };
    bins WkupHighSensitivityCalibInit                                 = { [ (('h40004278 - 'h40000000) >> 1) : ((('h40004278 - 'h40000000 + 'd92) >> 1) - 1) ] };
    bins McuRomCopyTxToRxCh37Dco                                      = { [ (('h400042d8 - 'h40000000) >> 1) : ((('h400042d8 - 'h40000000 + 'd62) >> 1) - 1) ] };
    bins McuRomCopyRxToTxCh37Dco                                      = { [ (('h40004318 - 'h40000000) >> 1) : ((('h40004318 - 'h40000000 + 'd62) >> 1) - 1) ] };
    bins SaveTxDcoForBleChannel                                       = { [ (('h40004358 - 'h40000000) >> 1) : ((('h40004358 - 'h40000000 + 'd232) >> 1) - 1) ] };
    bins RestoreTxDcoForBleChannel                                    = { [ (('h40004440 - 'h40000000) >> 1) : ((('h40004440 - 'h40000000 + 'd154) >> 1) - 1) ] };
    bins SetTxDcoForBleChannel                                        = { [ (('h400044e0 - 'h40000000) >> 1) : ((('h400044e0 - 'h40000000 + 'd94) >> 1) - 1) ] };
    bins GetTxDcoForBleChannel                                        = { [ (('h40004540 - 'h40000000) >> 1) : ((('h40004540 - 'h40000000 + 'd118) >> 1) - 1) ] };
    bins SetMinTxFreqForBleChannel                                    = { [ (('h400045b8 - 'h40000000) >> 1) : ((('h400045b8 - 'h40000000 + 'd118) >> 1) - 1) ] };
    bins SetMaxTxFreqForBleChannel                                    = { [ (('h40004630 - 'h40000000) >> 1) : ((('h40004630 - 'h40000000 + 'd94) >> 1) - 1) ] };
    bins DcoHop                                                       = { [ (('h40004690 - 'h40000000) >> 1) : ((('h40004690 - 'h40000000 + 'd432) >> 1) - 1) ] };
    bins DcoHopTxDcoEfine                                             = { [ (('h40004840 - 'h40000000) >> 1) : ((('h40004840 - 'h40000000 + 'd192) >> 1) - 1) ] };
    bins DcoHopTxDcoFine                                              = { [ (('h40004900 - 'h40000000) >> 1) : ((('h40004900 - 'h40000000 + 'd192) >> 1) - 1) ] };
    bins CalcEffEfine                                                 = { [ (('h400049c0 - 'h40000000) >> 1) : ((('h400049c0 - 'h40000000 + 'd172) >> 1) - 1) ] };
    bins FlowCopyAuxMeasureAndUnscaledToOvlMeasCtl                    = { [ (('h40004a70 - 'h40000000) >> 1) : ((('h40004a70 - 'h40000000 + 'd34) >> 1) - 1) ] };
    bins FlowSaveAuxMeasureAndUnscaledFromOvlMeasResult               = { [ (('h40004a98 - 'h40000000) >> 1) : ((('h40004a98 - 'h40000000 + 'd34) >> 1) - 1) ] };
    bins FlowCopyAuxMeasureToOvlMeasResult                            = { [ (('h40004ac0 - 'h40000000) >> 1) : ((('h40004ac0 - 'h40000000 + 'd14) >> 1) - 1) ] };
    bins EstimateAuxFreqFromAuxMeas                                   = { [ (('h40004ad0 - 'h40000000) >> 1) : ((('h40004ad0 - 'h40000000 + 'd20) >> 1) - 1) ] };
    bins CheckSwSideInfoFailOnChannel                                 = { [ (('h40004ae8 - 'h40000000) >> 1) : ((('h40004ae8 - 'h40000000 + 'd84) >> 1) - 1) ] };
    bins UpdateAuxMeasFromBleCh                                       = { [ (('h40004b40 - 'h40000000) >> 1) : ((('h40004b40 - 'h40000000 + 'd38) >> 1) - 1) ] };
    bins CheckSwSideInfoFail                                          = { [ (('h40004b68 - 'h40000000) >> 1) : ((('h40004b68 - 'h40000000 + 'd376) >> 1) - 1) ] };
    bins PrepareSecondDfMeas                                          = { [ (('h40004ce0 - 'h40000000) >> 1) : ((('h40004ce0 - 'h40000000 + 'd184) >> 1) - 1) ] };
    bins CalcDfandSprinklerStep                                       = { [ (('h40004d98 - 'h40000000) >> 1) : ((('h40004d98 - 'h40000000 + 'd336) >> 1) - 1) ] };
    bins McuRomDebugStuckMcuFunction                                  = { [ (('h40004ee8 - 'h40000000) >> 1) : ((('h40004ee8 - 'h40000000 + 'd54) >> 1) - 1) ] };
    bins DumpToDebugRam                                               = { [ (('h40004f20 - 'h40000000) >> 1) : ((('h40004f20 - 'h40000000 + 'd20) >> 1) - 1) ] };
    bins HwsJumpToSpecificRdr                                         = { [ (('h40004f38 - 'h40000000) >> 1) : ((('h40004f38 - 'h40000000 + 'd54) >> 1) - 1) ] };
    bins HwsJumpXRdrs                                                 = { [ (('h40004f70 - 'h40000000) >> 1) : ((('h40004f70 - 'h40000000 + 'd82) >> 1) - 1) ] };
    bins HwsNetJumpBack2Rdrs                                          = { [ (('h40004fc8 - 'h40000000) >> 1) : ((('h40004fc8 - 'h40000000 + 'd82) >> 1) - 1) ] };
    bins HwsNetJumpBack4Rdrs                                          = { [ (('h40005020 - 'h40000000) >> 1) : ((('h40005020 - 'h40000000 + 'd82) >> 1) - 1) ] };
    bins HwsNetJumpForward2Rdrs                                       = { [ (('h40005078 - 'h40000000) >> 1) : ((('h40005078 - 'h40000000 + 'd82) >> 1) - 1) ] };
    bins HwsNetJumpForward4Rdrs                                       = { [ (('h400050d0 - 'h40000000) >> 1) : ((('h400050d0 - 'h40000000 + 'd82) >> 1) - 1) ] };
    bins mcuRomDummyFunc                                              = { [ (('h40005128 - 'h40000000) >> 1) : ((('h40005128 - 'h40000000 + 'd46) >> 1) - 1) ] };
    bins McuRomWkupStateRoundRobinBleChannels                         = { [ (('h40005158 - 'h40000000) >> 1) : ((('h40005158 - 'h40000000 + 'd120) >> 1) - 1) ] };
    bins McuRomResetCalibParams                                       = { [ (('h400051d0 - 'h40000000) >> 1) : ((('h400051d0 - 'h40000000 + 'd100) >> 1) - 1) ] };
    bins StuckMCU                                                     = { [ (('h40005238 - 'h40000000) >> 1) : ((('h40005238 - 'h40000000 + 'd38) >> 1) - 1) ] };
    bins McuRomE4E4TestFunction                                       = { [ (('h40005260 - 'h40000000) >> 1) : ((('h40005260 - 'h40000000 + 'd38) >> 1) - 1) ] };
    bins McuRomFlowFSMPowerup                                         = { [ (('h40005288 - 'h40000000) >> 1) : ((('h40005288 - 'h40000000 + 'd430) >> 1) - 1) ] };
    bins McuRomResetLoVrefVbpAndLcAuxGnvmValues                       = { [ (('h40005438 - 'h40000000) >> 1) : ((('h40005438 - 'h40000000 + 'd32) >> 1) - 1) ] };
    bins McuRomSetEfineSteps                                          = { [ (('h40005458 - 'h40000000) >> 1) : ((('h40005458 - 'h40000000 + 'd30) >> 1) - 1) ] };
    bins McuRomSetParamsForFirstCycle                                 = { [ (('h40005478 - 'h40000000) >> 1) : ((('h40005478 - 'h40000000 + 'd2) >> 1) - 1) ] };
    bins McuRomRestoreParamsAfterFirstCycle                           = { [ (('h40005480 - 'h40000000) >> 1) : ((('h40005480 - 'h40000000 + 'd2) >> 1) - 1) ] };
    bins McuRomSetParamsForFirstPacket                                = { [ (('h40005488 - 'h40000000) >> 1) : ((('h40005488 - 'h40000000 + 'd28) >> 1) - 1) ] };
    bins McuRomRestoreParamsAfterFirstPacket                          = { [ (('h400054a8 - 'h40000000) >> 1) : ((('h400054a8 - 'h40000000 + 'd84) >> 1) - 1) ] };
    bins McuRomUpdateAuxMeasEstAndRxCalibUponNoTwoWU                  = { [ (('h40005500 - 'h40000000) >> 1) : ((('h40005500 - 'h40000000 + 'd94) >> 1) - 1) ] };
    bins McuRomTempSensingPowerUpConfig                               = { [ (('h40005560 - 'h40000000) >> 1) : ((('h40005560 - 'h40000000 + 'd104) >> 1) - 1) ] };
    bins McuRomAccTempSenseMeasInOvl                                  = { [ (('h400055c8 - 'h40000000) >> 1) : ((('h400055c8 - 'h40000000 + 'd64) >> 1) - 1) ] };
    bins McuRomTempChangeEvent                                        = { [ (('h40005608 - 'h40000000) >> 1) : ((('h40005608 - 'h40000000 + 'd254) >> 1) - 1) ] };
    bins McuRomCalcTempFromSensorFsm                                  = { [ (('h40005708 - 'h40000000) >> 1) : ((('h40005708 - 'h40000000 + 'd394) >> 1) - 1) ] };
    bins McuRomTempComp                                               = { [ (('h40005898 - 'h40000000) >> 1) : ((('h40005898 - 'h40000000 + 'd100) >> 1) - 1) ] };
    bins McuRomSetAdbDoneDelayUponFirstTempComp                       = { [ (('h40005900 - 'h40000000) >> 1) : ((('h40005900 - 'h40000000 + 'd42) >> 1) - 1) ] };
    bins McuRomAdbDoneDelayTempComp                                   = { [ (('h40005930 - 'h40000000) >> 1) : ((('h40005930 - 'h40000000 + 'd156) >> 1) - 1) ] };
    bins McuRomRcSensingPowerUpConfig                                 = { [ (('h400059d0 - 'h40000000) >> 1) : ((('h400059d0 - 'h40000000 + 'd62) >> 1) - 1) ] };
    bins McuRomRcSensingFsm                                           = { [ (('h40005a10 - 'h40000000) >> 1) : ((('h40005a10 - 'h40000000 + 'd478) >> 1) - 1) ] };
    bins McuRomRoundRobinRCSensorConfig                               = { [ (('h40005bf0 - 'h40000000) >> 1) : ((('h40005bf0 - 'h40000000 + 'd88) >> 1) - 1) ] };
    bins McuRomTamperSensing                                          = { [ (('h40005c48 - 'h40000000) >> 1) : ((('h40005c48 - 'h40000000 + 'd100) >> 1) - 1) ] };
    bins McuRomCalcNumEnvDetsCyclesForBle5                            = { [ (('h40005cb0 - 'h40000000) >> 1) : ((('h40005cb0 - 'h40000000 + 'd222) >> 1) - 1) ] };
    bins McuRomRestoreFromFastEnvdetClk                               = { [ (('h40005d90 - 'h40000000) >> 1) : ((('h40005d90 - 'h40000000 + 'd156) >> 1) - 1) ] };
    bins McuRomLoVrefVbpCalibCleFsm                                   = { [ (('h40005e30 - 'h40000000) >> 1) : ((('h40005e30 - 'h40000000 + 'd1162) >> 1) - 1) ] };
    bins McuRomLoVrefVbpCalibCleFsmWithCh39                           = { [ (('h400062c0 - 'h40000000) >> 1) : ((('h400062c0 - 'h40000000 + 'd834) >> 1) - 1) ] };
    bins McuRomLoVrefVbpCalibCleFsmE2                                 = { [ (('h40006608 - 'h40000000) >> 1) : ((('h40006608 - 'h40000000 + 'd648) >> 1) - 1) ] };
    bins McuRomLoVrefVbpCalibFsm                                      = { [ (('h40006890 - 'h40000000) >> 1) : ((('h40006890 - 'h40000000 + 'd860) >> 1) - 1) ] };
    bins McuRomForceVrefVbpWithoutCalib                               = { [ (('h40006bf0 - 'h40000000) >> 1) : ((('h40006bf0 - 'h40000000 + 'd74) >> 1) - 1) ] };
    bins McuRomLcAuxCalibCleFsm                                       = { [ (('h40006c40 - 'h40000000) >> 1) : ((('h40006c40 - 'h40000000 + 'd578) >> 1) - 1) ] };
    bins McuRomLcAuxCalibFsm                                          = { [ (('h40006e88 - 'h40000000) >> 1) : ((('h40006e88 - 'h40000000 + 'd554) >> 1) - 1) ] };
    bins McuRomDfAndSprinklerStepCalibFsm                             = { [ (('h400070b8 - 'h40000000) >> 1) : ((('h400070b8 - 'h40000000 + 'd914) >> 1) - 1) ] };
    bins McuRomDfConfigBetweenConsecMeas                              = { [ (('h40007450 - 'h40000000) >> 1) : ((('h40007450 - 'h40000000 + 'd112) >> 1) - 1) ] };
    bins McuRomLoTxRxCalibPreProcessing                               = { [ (('h400074c0 - 'h40000000) >> 1) : ((('h400074c0 - 'h40000000 + 'd122) >> 1) - 1) ] };
    bins McuRomLoTxRxCalibPostProcessing                              = { [ (('h40007540 - 'h40000000) >> 1) : ((('h40007540 - 'h40000000 + 'd312) >> 1) - 1) ] };
    bins McuRomLoCalibFsm                                             = { [ (('h40007678 - 'h40000000) >> 1) : ((('h40007678 - 'h40000000 + 'd864) >> 1) - 1) ] };
    bins McuRomLoCalibFsmE2                                           = { [ (('h400079d8 - 'h40000000) >> 1) : ((('h400079d8 - 'h40000000 + 'd558) >> 1) - 1) ] };
    bins McuRomCopyCalibRsltCoarseToHrr                               = { [ (('h40007c08 - 'h40000000) >> 1) : ((('h40007c08 - 'h40000000 + 'd92) >> 1) - 1) ] };
    bins McuRomUpdatePacketDataForTestMode                            = { [ (('h40007c68 - 'h40000000) >> 1) : ((('h40007c68 - 'h40000000 + 'd2) >> 1) - 1) ] };
    bins McuRomPostPacketPreparation                                  = { [ (('h40007c70 - 'h40000000) >> 1) : ((('h40007c70 - 'h40000000 + 'd200) >> 1) - 1) ] };
    bins McuRomSaveHalfMic                                            = { [ (('h40007d38 - 'h40000000) >> 1) : ((('h40007d38 - 'h40000000 + 'd28) >> 1) - 1) ] };
    bins McuRomCombineTwoMics                                         = { [ (('h40007d58 - 'h40000000) >> 1) : ((('h40007d58 - 'h40000000 + 'd48) >> 1) - 1) ] };
    bins McuRomUpdateNonceForPacketType                               = { [ (('h40007d88 - 'h40000000) >> 1) : ((('h40007d88 - 'h40000000 + 'd30) >> 1) - 1) ] };
    bins McuRomUpdatePacketTypeInGroupId                              = { [ (('h40007da8 - 'h40000000) >> 1) : ((('h40007da8 - 'h40000000 + 'd30) >> 1) - 1) ] };
    bins McuRomUpdatePacketData                                       = { [ (('h40007dc8 - 'h40000000) >> 1) : ((('h40007dc8 - 'h40000000 + 'd776) >> 1) - 1) ] };
    bins McuRomUpdatePacketDataForMiniRx                              = { [ (('h400080d0 - 'h40000000) >> 1) : ((('h400080d0 - 'h40000000 + 'd122) >> 1) - 1) ] };
    bins McuRomTxSprinkler                                            = { [ (('h40008150 - 'h40000000) >> 1) : ((('h40008150 - 'h40000000 + 'd766) >> 1) - 1) ] };
    bins McuRomSetRegsForExtendedPacket                               = { [ (('h40008450 - 'h40000000) >> 1) : ((('h40008450 - 'h40000000 + 'd70) >> 1) - 1) ] };
    bins McuRomTxBle5SetParams                                        = { [ (('h40008498 - 'h40000000) >> 1) : ((('h40008498 - 'h40000000 + 'd318) >> 1) - 1) ] };
    bins McuRomTxBle5SetWkupParams                                    = { [ (('h400085d8 - 'h40000000) >> 1) : ((('h400085d8 - 'h40000000 + 'd216) >> 1) - 1) ] };
    bins McuRomTxBle5SetRadioParams                                   = { [ (('h400086b0 - 'h40000000) >> 1) : ((('h400086b0 - 'h40000000 + 'd108) >> 1) - 1) ] };
    bins McuRomTxBle5RestoreParams                                    = { [ (('h40008720 - 'h40000000) >> 1) : ((('h40008720 - 'h40000000 + 'd104) >> 1) - 1) ] };
    bins McuRomBle5CheckSoftAwdtInd                                   = { [ (('h40008788 - 'h40000000) >> 1) : ((('h40008788 - 'h40000000 + 'd116) >> 1) - 1) ] };
    bins McuRomSetAwdtForBle5DataPacket                               = { [ (('h40008800 - 'h40000000) >> 1) : ((('h40008800 - 'h40000000 + 'd42) >> 1) - 1) ] };
    bins McuRomFlowManagerDebugUpdateMaskUponCycleBegin               = { [ (('h40008830 - 'h40000000) >> 1) : ((('h40008830 - 'h40000000 + 'd74) >> 1) - 1) ] };
    bins McuRomFlowManagerDisableJumpForGivenState                    = { [ (('h40008880 - 'h40000000) >> 1) : ((('h40008880 - 'h40000000 + 'd78) >> 1) - 1) ] };
    bins McuRomPreLoProximityMeas                                     = { [ (('h400088d0 - 'h40000000) >> 1) : ((('h400088d0 - 'h40000000 + 'd152) >> 1) - 1) ] };
    bins McuRomPostLoProximityMeas                                    = { [ (('h40008968 - 'h40000000) >> 1) : ((('h40008968 - 'h40000000 + 'd266) >> 1) - 1) ] };
    bins McuRomLoProximityCheckScanDcoMode                            = { [ (('h40008a78 - 'h40000000) >> 1) : ((('h40008a78 - 'h40000000 + 'd88) >> 1) - 1) ] };
    bins McuRomPostLoProximityMeasForDcoScan                          = { [ (('h40008ad0 - 'h40000000) >> 1) : ((('h40008ad0 - 'h40000000 + 'd78) >> 1) - 1) ] };
    bins McuRomCloseWkup                                              = { [ (('h40008b20 - 'h40000000) >> 1) : ((('h40008b20 - 'h40000000 + 'd26) >> 1) - 1) ] };
    bins McuRomSetLoDcoCoarseForWkup                                  = { [ (('h40008b40 - 'h40000000) >> 1) : ((('h40008b40 - 'h40000000 + 'd206) >> 1) - 1) ] };
    bins McuRomRestoreLoDcoCoarseAfterWkup                            = { [ (('h40008c10 - 'h40000000) >> 1) : ((('h40008c10 - 'h40000000 + 'd54) >> 1) - 1) ] };
    bins McuRomPrepareForWkupCh37Event                                = { [ (('h40008c48 - 'h40000000) >> 1) : ((('h40008c48 - 'h40000000 + 'd12) >> 1) - 1) ] };
    bins McuRomPrepareForWkupCh38Event                                = { [ (('h40008c58 - 'h40000000) >> 1) : ((('h40008c58 - 'h40000000 + 'd12) >> 1) - 1) ] };
    bins McuRomPrepareForWkupCh39Event                                = { [ (('h40008c68 - 'h40000000) >> 1) : ((('h40008c68 - 'h40000000 + 'd12) >> 1) - 1) ] };
    bins McuRomSaveChargingTime                                       = { [ (('h40008c78 - 'h40000000) >> 1) : ((('h40008c78 - 'h40000000 + 'd56) >> 1) - 1) ] };
    bins McuRomSaveEAWKUPTimers                                       = { [ (('h40008cb0 - 'h40000000) >> 1) : ((('h40008cb0 - 'h40000000 + 'd38) >> 1) - 1) ] };
    bins McuRomSetParamsForCcaSequence                                = { [ (('h40008cd8 - 'h40000000) >> 1) : ((('h40008cd8 - 'h40000000 + 'd116) >> 1) - 1) ] };
    bins McuRomEnvdetClkConfigPostMeas                                = { [ (('h40008d50 - 'h40000000) >> 1) : ((('h40008d50 - 'h40000000 + 'd78) >> 1) - 1) ] };
    bins McuRomSetParamsForWkupSequence                               = { [ (('h40008da0 - 'h40000000) >> 1) : ((('h40008da0 - 'h40000000 + 'd122) >> 1) - 1) ] };
    bins McuRomSystemClksMeasFsm                                      = { [ (('h40008e20 - 'h40000000) >> 1) : ((('h40008e20 - 'h40000000 + 'd520) >> 1) - 1) ] };
    bins McuRomSetFastEnvdetClk                                       = { [ (('h40009028 - 'h40000000) >> 1) : ((('h40009028 - 'h40000000 + 'd106) >> 1) - 1) ] };
    bins McuRomEnvdetClkConfigPreMeas                                 = { [ (('h40009098 - 'h40000000) >> 1) : ((('h40009098 - 'h40000000 + 'd126) >> 1) - 1) ] };
    bins McuRomWkupCalibCleFsm                                        = { [ (('h40009118 - 'h40000000) >> 1) : ((('h40009118 - 'h40000000 + 'd626) >> 1) - 1) ] };
    bins McuRomWkupLowSensitivityCalibFsm                             = { [ (('h40009390 - 'h40000000) >> 1) : ((('h40009390 - 'h40000000 + 'd428) >> 1) - 1) ] };
    bins McuRomWkupHighSensitivityCalibFsm                            = { [ (('h40009540 - 'h40000000) >> 1) : ((('h40009540 - 'h40000000 + 'd592) >> 1) - 1) ] };
    bins McuRomWkupCalibFsm                                           = { [ (('h40009790 - 'h40000000) >> 1) : ((('h40009790 - 'h40000000 + 'd30) >> 1) - 1) ] };
    bins SetBasicFlowWUParams                                         = { [ (('h400097b0 - 'h40000000) >> 1) : ((('h400097b0 - 'h40000000 + 'd64) >> 1) - 1) ] };
    bins FlowDCOSetCH37                                               = { [ (('h400097f0 - 'h40000000) >> 1) : ((('h400097f0 - 'h40000000 + 'd10) >> 1) - 1) ] };
    bins FlowDCOSetCH38                                               = { [ (('h40009800 - 'h40000000) >> 1) : ((('h40009800 - 'h40000000 + 'd12) >> 1) - 1) ] };
    bins FlowDCOSetCH39                                               = { [ (('h40009810 - 'h40000000) >> 1) : ((('h40009810 - 'h40000000 + 'd12) >> 1) - 1) ] };
    bins McuRomChannelHopping                                         = { [ (('h40009820 - 'h40000000) >> 1) : ((('h40009820 - 'h40000000 + 'd42) >> 1) - 1) ] };
    bins PerformSwAlphaFiltering                                      = { [ (('h40009850 - 'h40000000) >> 1) : ((('h40009850 - 'h40000000 + 'd66) >> 1) - 1) ] };
    bins McuRomClearSwspad31                                          = { [ (('h40009898 - 'h40000000) >> 1) : ((('h40009898 - 'h40000000 + 'd10) >> 1) - 1) ] };
    bins FlowJump                                                     = { [ (('h400098a8 - 'h40000000) >> 1) : ((('h400098a8 - 'h40000000 + 'd20) >> 1) - 1) ] };
    bins McuRomEvaluateSystemTime                                     = { [ (('h400098c0 - 'h40000000) >> 1) : ((('h400098c0 - 'h40000000 + 'd218) >> 1) - 1) ] };
    bins McuRomFlowManagerFsm                                         = { [ (('h400099a0 - 'h40000000) >> 1) : ((('h400099a0 - 'h40000000 + 'd1850) >> 1) - 1) ] };
    bins McuRomUpdateAdvaFromNonce                                    = { [ (('h4000a0e0 - 'h40000000) >> 1) : ((('h4000a0e0 - 'h40000000 + 'd32) >> 1) - 1) ] };
    bins McuRomSetTxRxParamsForAuxMeas                                = { [ (('h4000a100 - 'h40000000) >> 1) : ((('h4000a100 - 'h40000000 + 'd94) >> 1) - 1) ] };
    bins McuRomRestoreTxRxParamsAfterAuxMeas                          = { [ (('h4000a160 - 'h40000000) >> 1) : ((('h4000a160 - 'h40000000 + 'd64) >> 1) - 1) ] };
    bins McuRomAuxMeasFsm                                             = { [ (('h4000a1a0 - 'h40000000) >> 1) : ((('h4000a1a0 - 'h40000000 + 'd622) >> 1) - 1) ] };
    bins McuCopyCalibRsltCoarseToHrr                                  = { [ (('h4000a410 - 'h40000000) >> 1) : ((('h4000a410 - 'h40000000 + 'd92) >> 1) - 1) ] };
    bins McuBasicFlowCheckTxTimeSprinkler                             = { [ (('h4000a470 - 'h40000000) >> 1) : ((('h4000a470 - 'h40000000 + 'd70) >> 1) - 1) ] };
    bins McuBasicFlowCheckIfSymCalibEn                                = { [ (('h4000a4b8 - 'h40000000) >> 1) : ((('h4000a4b8 - 'h40000000 + 'd26) >> 1) - 1) ] };
    bins McuBasicFlowChoseSymForPgx                                   = { [ (('h4000a4d8 - 'h40000000) >> 1) : ((('h4000a4d8 - 'h40000000 + 'd26) >> 1) - 1) ] };
    bins McuRomBasicFlowUpdateAuxMeas                                 = { [ (('h4000a4f8 - 'h40000000) >> 1) : ((('h4000a4f8 - 'h40000000 + 'd48) >> 1) - 1) ] };
    bins McuBasicFlowSetLoDiv2Sym                                     = { [ (('h4000a528 - 'h40000000) >> 1) : ((('h4000a528 - 'h40000000 + 'd62) >> 1) - 1) ] };
    bins McuRomBasicFlowBuildPacket                                   = { [ (('h4000a568 - 'h40000000) >> 1) : ((('h4000a568 - 'h40000000 + 'd168) >> 1) - 1) ] };
    bins McuRomBasicFlowSetRoundRobin                                 = { [ (('h4000a610 - 'h40000000) >> 1) : ((('h4000a610 - 'h40000000 + 'd40) >> 1) - 1) ] };
    bins McuRomBasicFlowCheck2WU                                      = { [ (('h4000a638 - 'h40000000) >> 1) : ((('h4000a638 - 'h40000000 + 'd152) >> 1) - 1) ] };
    bins McuRomSetWkupParamsPreRx                                     = { [ (('h4000a6d0 - 'h40000000) >> 1) : ((('h4000a6d0 - 'h40000000 + 'd38) >> 1) - 1) ] };
    bins McuRomMiniRxFSM                                              = { [ (('h4000a6f8 - 'h40000000) >> 1) : ((('h4000a6f8 - 'h40000000 + 'd472) >> 1) - 1) ] };
    bins McuRomMiniRxStoreWkupParams                                  = { [ (('h4000a8d0 - 'h40000000) >> 1) : ((('h4000a8d0 - 'h40000000 + 'd198) >> 1) - 1) ] };
    bins McuRomMiniRxRestoreWkupParams                                = { [ (('h4000a998 - 'h40000000) >> 1) : ((('h4000a998 - 'h40000000 + 'd104) >> 1) - 1) ] };
    bins McuRomMiniRxCheckDone                                        = { [ (('h4000aa00 - 'h40000000) >> 1) : ((('h4000aa00 - 'h40000000 + 'd284) >> 1) - 1) ] };
    bins McuRomMiniRxDebugPowerGearConfig                             = { [ (('h4000ab20 - 'h40000000) >> 1) : ((('h4000ab20 - 'h40000000 + 'd28) >> 1) - 1) ] };
    bins McuRomSetEnterTestModeParams                                 = { [ (('h4000ab40 - 'h40000000) >> 1) : ((('h4000ab40 - 'h40000000 + 'd94) >> 1) - 1) ] };
    bins McuRomTestModeResetTO                                        = { [ (('h4000aba0 - 'h40000000) >> 1) : ((('h4000aba0 - 'h40000000 + 'd30) >> 1) - 1) ] };
    bins McuRomCheckTestModeTimeOut                                   = { [ (('h4000abc0 - 'h40000000) >> 1) : ((('h4000abc0 - 'h40000000 + 'd56) >> 1) - 1) ] };
    bins McuRomCheckMeasuredValueTestMode                             = { [ (('h4000abf8 - 'h40000000) >> 1) : ((('h4000abf8 - 'h40000000 + 'd260) >> 1) - 1) ] };
    bins McuRomTestModeCheckWUStateReached                            = { [ (('h4000ad00 - 'h40000000) >> 1) : ((('h4000ad00 - 'h40000000 + 'd28) >> 1) - 1) ] };
    bins McuRomSetCwScalerForTestMode                                 = { [ (('h4000ad20 - 'h40000000) >> 1) : ((('h4000ad20 - 'h40000000 + 'd48) >> 1) - 1) ] };
    bins McuRomUpdateTestModePacketAndSetLoDiv2Sym                    = { [ (('h4000ad50 - 'h40000000) >> 1) : ((('h4000ad50 - 'h40000000 + 'd204) >> 1) - 1) ] };
    bins McuRomRestoreParamsAfterTestmode                             = { [ (('h4000ae20 - 'h40000000) >> 1) : ((('h4000ae20 - 'h40000000 + 'd86) >> 1) - 1) ] };
    bins McuRomCheckSprinklerTestmode                                 = { [ (('h4000ae78 - 'h40000000) >> 1) : ((('h4000ae78 - 'h40000000 + 'd40) >> 1) - 1) ] };
    bins McuRomDebugSetMiniRxStateInLoProx                            = { [ (('h4000aea0 - 'h40000000) >> 1) : ((('h4000aea0 - 'h40000000 + 'd20) >> 1) - 1) ] };
    bins McuRomSetTestUpdateSprinklerAndUID                           = { [ (('h4000aeb8 - 'h40000000) >> 1) : ((('h4000aeb8 - 'h40000000 + 'd44) >> 1) - 1) ] };
    bins McuRomTestModeCheckBeaconLengthBelowTH                       = { [ (('h4000aee8 - 'h40000000) >> 1) : ((('h4000aee8 - 'h40000000 + 'd130) >> 1) - 1) ] };
    bins McuRomTestModeEstimateFrequencyDelta                         = { [ (('h4000af70 - 'h40000000) >> 1) : ((('h4000af70 - 'h40000000 + 'd50) >> 1) - 1) ] };
    bins McuRomTestModeCheckIfEnterFrequency                          = { [ (('h4000afa8 - 'h40000000) >> 1) : ((('h4000afa8 - 'h40000000 + 'd96) >> 1) - 1) ] };
    bins McuRomTestModeValidateEnterFrequencyDelta                    = { [ (('h4000b008 - 'h40000000) >> 1) : ((('h4000b008 - 'h40000000 + 'd86) >> 1) - 1) ] };
    bins McuRomTestModeCopyChannelYValToSWSPAD                        = { [ (('h4000b060 - 'h40000000) >> 1) : ((('h4000b060 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins McuRomHarvFlowCounter                                        = { [ (('h4000b0a0 - 'h40000000) >> 1) : ((('h4000b0a0 - 'h40000000 + 'd56) >> 1) - 1) ] };
    bins McuRomAddBitToMask                                           = { [ (('h4000b0d8 - 'h40000000) >> 1) : ((('h4000b0d8 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins McuRomJump2IfNotFirstCycle                                   = { [ (('h4000b118 - 'h40000000) >> 1) : ((('h4000b118 - 'h40000000 + 'd26) >> 1) - 1) ] };
    bins FlowInit_UID                                                 = { [ (('h4000b138 - 'h40000000) >> 1) : ((('h4000b138 - 'h40000000 + 'd18) >> 1) - 1) ] };
    bins McuRomInitSocClock                                           = { [ (('h4000b150 - 'h40000000) >> 1) : ((('h4000b150 - 'h40000000 + 'd2) >> 1) - 1) ] };
    bins McuRomSOCCalibration                                         = { [ (('h4000b158 - 'h40000000) >> 1) : ((('h4000b158 - 'h40000000 + 'd432) >> 1) - 1) ] };
    bins McuRomMeasureFreq                                            = { [ (('h4000b308 - 'h40000000) >> 1) : ((('h4000b308 - 'h40000000 + 'd274) >> 1) - 1) ] };
    bins McuRomBinarySearchFMU                                        = { [ (('h4000b41c - 'h40000000) >> 1) : ((('h4000b41c - 'h40000000 + 'd714) >> 1) - 1) ] };
    bins McuRomAfterBinarySearchControl                               = { [ (('h4000b6e8 - 'h40000000) >> 1) : ((('h4000b6e8 - 'h40000000 + 'd186) >> 1) - 1) ] };
    bins McuRomRTCCalibrationStore                                    = { [ (('h4000b7a4 - 'h40000000) >> 1) : ((('h4000b7a4 - 'h40000000 + 'd176) >> 1) - 1) ] };
    bins McuRomRTCCalibration                                         = { [ (('h4000b858 - 'h40000000) >> 1) : ((('h4000b858 - 'h40000000 + 'd554) >> 1) - 1) ] };
    bins McuRomWURXCalibration                                        = { [ (('h4000ba84 - 'h40000000) >> 1) : ((('h4000ba84 - 'h40000000 + 'd476) >> 1) - 1) ] };
    bins McuRomActiveCalibration                                      = { [ (('h4000bc60 - 'h40000000) >> 1) : ((('h4000bc60 - 'h40000000 + 'd336) >> 1) - 1) ] };
    bins McuRomRunFMU                                                 = { [ (('h4000bdb0 - 'h40000000) >> 1) : ((('h4000bdb0 - 'h40000000 + 'd140) >> 1) - 1) ] };
    bins McuRomFmuCmd                                                 = { [ (('h4000be3c - 'h40000000) >> 1) : ((('h4000be3c - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins McuRomOtpBlockCompare                                        = { [ (('h4000be4c - 'h40000000) >> 1) : ((('h4000be4c - 'h40000000 + 'd92) >> 1) - 1) ] };
    bins McuRomCalcBer                                                = { [ (('h4000bea8 - 'h40000000) >> 1) : ((('h4000bea8 - 'h40000000 + 'd30) >> 1) - 1) ] };
    bins WriteToAddr                                                  = { [ (('h4000bec8 - 'h40000000) >> 1) : ((('h4000bec8 - 'h40000000 + 'd18) >> 1) - 1) ] };
    bins GetFromAddr                                                  = { [ (('h4000bedc - 'h40000000) >> 1) : ((('h4000bedc - 'h40000000 + 'd10) >> 1) - 1) ] };
    bins SetRadioInitTableAddress                                     = { [ (('h4000bee8 - 'h40000000) >> 1) : ((('h4000bee8 - 'h40000000 + 'd42) >> 1) - 1) ] };
    bins CopyRadioModeRegister                                        = { [ (('h4000bf14 - 'h40000000) >> 1) : ((('h4000bf14 - 'h40000000 + 'd14) >> 1) - 1) ] };
    bins EnableExtAndSwEvents                                         = { [ (('h4000bf24 - 'h40000000) >> 1) : ((('h4000bf24 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins setDelay                                                     = { [ (('h4000bf34 - 'h40000000) >> 1) : ((('h4000bf34 - 'h40000000 + 'd40) >> 1) - 1) ] };
    bins WaitForDelay                                                 = { [ (('h4000bf5c - 'h40000000) >> 1) : ((('h4000bf5c - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins WaitForSysEventWithTimeOut                                   = { [ (('h4000bf98 - 'h40000000) >> 1) : ((('h4000bf98 - 'h40000000 + 'd104) >> 1) - 1) ] };
    bins McuRomHwsJumpXRdrs_RelativeToFunc                            = { [ (('h4000c000 - 'h40000000) >> 1) : ((('h4000c000 - 'h40000000 + 'd80) >> 1) - 1) ] };
    bins ExceptionHandlerDefault                                      = { [ (('h4000cb00 - 'h40000000) >> 1) : ((('h4000cb00 - 'h40000000 + 'd8) >> 1) - 1) ] };
    bins abs                                                          = { [ (('h4000cb0c - 'h40000000) >> 1) : ((('h4000cb0c - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins div                                                          = { [ (('h4000cb1c - 'h40000000) >> 1) : ((('h4000cb1c - 'h40000000 + 'd72) >> 1) - 1) ] };
    bins memchr                                                       = { [ (('h4000cb64 - 'h40000000) >> 1) : ((('h4000cb64 - 'h40000000 + 'd200) >> 1) - 1) ] };
    bins memcmp                                                       = { [ (('h4000cc2c - 'h40000000) >> 1) : ((('h4000cc2c - 'h40000000 + 'd120) >> 1) - 1) ] };
    bins memcpy                                                       = { [ (('h4000cca4 - 'h40000000) >> 1) : ((('h4000cca4 - 'h40000000 + 'd428) >> 1) - 1) ] };
    bins memmove                                                      = { [ (('h4000ce50 - 'h40000000) >> 1) : ((('h4000ce50 - 'h40000000 + 'd332) >> 1) - 1) ] };
    bins memset                                                       = { [ (('h4000cf9c - 'h40000000) >> 1) : ((('h4000cf9c - 'h40000000 + 'd220) >> 1) - 1) ] };
    bins srand                                                        = { [ (('h4000d078 - 'h40000000) >> 1) : ((('h4000d078 - 'h40000000 + 'd20) >> 1) - 1) ] };
    bins rand                                                         = { [ (('h4000d08c - 'h40000000) >> 1) : ((('h4000d08c - 'h40000000 + 'd88) >> 1) - 1) ] };
    bins McuDramAdcCompGo                                             = { [ (('h40010000 - 'h40000000) >> 1) : ((('h40010000 - 'h40000000 + 'd106) >> 1) - 1) ] };
    bins McuDramInitSrrForVtest                                       = { [ (('h40010000 - 'h40000000) >> 1) : ((('h40010000 - 'h40000000 + 'd34) >> 1) - 1) ] };
    bins McuDramSetTempSensDemLenDemCtl                               = { [ (('h40010000 - 'h40000000) >> 1) : ((('h40010000 - 'h40000000 + 'd46) >> 1) - 1) ] };
    bins McuDramSystemClocksCalibration                               = { [ (('h40010000 - 'h40000000) >> 1) : ((('h40010000 - 'h40000000 + 'd438) >> 1) - 1) ] };
    bins McuDramSystemClocksCharacterization                          = { [ (('h40010000 - 'h40000000) >> 1) : ((('h40010000 - 'h40000000 + 'd160) >> 1) - 1) ] };
    bins McuDramWkupDiv2Verify                                        = { [ (('h40010000 - 'h40000000) >> 1) : ((('h40010000 - 'h40000000 + 'd320) >> 1) - 1) ] };
    bins McuDramWsVstartCalib                                         = { [ (('h40010000 - 'h40000000) >> 1) : ((('h40010000 - 'h40000000 + 'd274) >> 1) - 1) ] };
    bins MCU_Exception_Handler                                        = { [ (('h40010000 - 'h40000000) >> 1) : ((('h40010000 - 'h40000000 + 'd44) >> 1) - 1) ] };
    bins McuDramValidateRetValuesAfterPoff                            = { [ (('h40010024 - 'h40000000) >> 1) : ((('h40010024 - 'h40000000 + 'd180) >> 1) - 1) ] };
    bins CheckInitial_AuxWU                                           = { [ (('h40010030 - 'h40000000) >> 1) : ((('h40010030 - 'h40000000 + 'd32) >> 1) - 1) ] };
    bins McuDramSetDem                                                = { [ (('h40010030 - 'h40000000) >> 1) : ((('h40010030 - 'h40000000 + 'd120) >> 1) - 1) ] };
    bins MCU_Set_WU_Configuration                                     = { [ (('h40010050 - 'h40000000) >> 1) : ((('h40010050 - 'h40000000 + 'd120) >> 1) - 1) ] };
    bins McuDramAdcCompCalc                                           = { [ (('h40010070 - 'h40000000) >> 1) : ((('h40010070 - 'h40000000 + 'd84) >> 1) - 1) ] };
    bins McuDramRTCChar                                               = { [ (('h400100a0 - 'h40000000) >> 1) : ((('h400100a0 - 'h40000000 + 'd386) >> 1) - 1) ] };
    bins McuDramCTATCalibrationFSM                                    = { [ (('h400100a8 - 'h40000000) >> 1) : ((('h400100a8 - 'h40000000 + 'd448) >> 1) - 1) ] };
    bins McuDramAdcCompCalcWrapper                                    = { [ (('h400100c8 - 'h40000000) >> 1) : ((('h400100c8 - 'h40000000 + 'd232) >> 1) - 1) ] };
    bins MCU_Set_WU                                                   = { [ (('h400100c8 - 'h40000000) >> 1) : ((('h400100c8 - 'h40000000 + 'd80) >> 1) - 1) ] };
    bins McuDramVerifyOtpEndlessRead                                  = { [ (('h400100d8 - 'h40000000) >> 1) : ((('h400100d8 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins McuSetParamsForSymMeasLc                                     = { [ (('h400100e8 - 'h40000000) >> 1) : ((('h400100e8 - 'h40000000 + 'd122) >> 1) - 1) ] };
    bins McuDramVstartVerif                                           = { [ (('h40010114 - 'h40000000) >> 1) : ((('h40010114 - 'h40000000 + 'd20) >> 1) - 1) ] };
    bins MCU_Set_CCA                                                  = { [ (('h40010118 - 'h40000000) >> 1) : ((('h40010118 - 'h40000000 + 'd26) >> 1) - 1) ] };
    bins McuDramVstartStore                                           = { [ (('h40010128 - 'h40000000) >> 1) : ((('h40010128 - 'h40000000 + 'd144) >> 1) - 1) ] };
    bins McuDramTempStaticCompFix                                     = { [ (('h40010134 - 'h40000000) >> 1) : ((('h40010134 - 'h40000000 + 'd130) >> 1) - 1) ] };
    bins McuSetParamsForLcCalibSym                                    = { [ (('h40010164 - 'h40000000) >> 1) : ((('h40010164 - 'h40000000 + 'd148) >> 1) - 1) ] };
    bins McuDramVddAdbCalib                                           = { [ (('h400101b0 - 'h40000000) >> 1) : ((('h400101b0 - 'h40000000 + 'd62) >> 1) - 1) ] };
    bins McuDramCalcTdcAndSetTrim                                     = { [ (('h400101b8 - 'h40000000) >> 1) : ((('h400101b8 - 'h40000000 + 'd974) >> 1) - 1) ] };
    bins McuDramInitRcSenseCalib                                      = { [ (('h400101b8 - 'h40000000) >> 1) : ((('h400101b8 - 'h40000000 + 'd26) >> 1) - 1) ] };
    bins McuDramSimpleDmaCommon                                       = { [ (('h400101b8 - 'h40000000) >> 1) : ((('h400101b8 - 'h40000000 + 'd42) >> 1) - 1) ] };
    bins McuDramRcSenseInit                                           = { [ (('h400101d4 - 'h40000000) >> 1) : ((('h400101d4 - 'h40000000 + 'd66) >> 1) - 1) ] };
    bins McuDramVddDigCalib                                           = { [ (('h400101f0 - 'h40000000) >> 1) : ((('h400101f0 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins McuNvmCopyAuxMeasToIsp                                       = { [ (('h400101f8 - 'h40000000) >> 1) : ((('h400101f8 - 'h40000000 + 'd80) >> 1) - 1) ] };
    bins McuDramRcSenseCheckResult                                    = { [ (('h40010218 - 'h40000000) >> 1) : ((('h40010218 - 'h40000000 + 'd288) >> 1) - 1) ] };
    bins McuDramSystemClocksCharacterizationRtc                       = { [ (('h40010222 - 'h40000000) >> 1) : ((('h40010222 - 'h40000000 + 'd74) >> 1) - 1) ] };
    bins McuDramVddSym600Calib                                        = { [ (('h40010230 - 'h40000000) >> 1) : ((('h40010230 - 'h40000000 + 'd56) >> 1) - 1) ] };
    bins McuNvmCopySymCalibResultsToIsp                               = { [ (('h40010248 - 'h40000000) >> 1) : ((('h40010248 - 'h40000000 + 'd178) >> 1) - 1) ] };
    bins McuDramAdjustJumpForCtatCalibSrrFlow                         = { [ (('h40010268 - 'h40000000) >> 1) : ((('h40010268 - 'h40000000 + 'd32) >> 1) - 1) ] };
    bins McuDramVddSym750Calib                                        = { [ (('h40010268 - 'h40000000) >> 1) : ((('h40010268 - 'h40000000 + 'd56) >> 1) - 1) ] };
    bins McuDramCalcCtrlChar                                          = { [ (('h4001026c - 'h40000000) >> 1) : ((('h4001026c - 'h40000000 + 'd88) >> 1) - 1) ] };
    bins McuDramVddCBias525Calib                                      = { [ (('h400102a0 - 'h40000000) >> 1) : ((('h400102a0 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins McuDramWURXCharacterization                                  = { [ (('h400102c4 - 'h40000000) >> 1) : ((('h400102c4 - 'h40000000 + 'd316) >> 1) - 1) ] };
    bins McuDramVddCBias175Calib                                      = { [ (('h400102e0 - 'h40000000) >> 1) : ((('h400102e0 - 'h40000000 + 'd82) >> 1) - 1) ] };
    bins McuDramLcAuxIdacCalibStore                                   = { [ (('h400102fc - 'h40000000) >> 1) : ((('h400102fc - 'h40000000 + 'd22) >> 1) - 1) ] };
    bins McuDramWkUpBbamp                                             = { [ (('h40010314 - 'h40000000) >> 1) : ((('h40010314 - 'h40000000 + 'd32) >> 1) - 1) ] };
    bins McuDramWkUpVerif                                             = { [ (('h40010334 - 'h40000000) >> 1) : ((('h40010334 - 'h40000000 + 'd30) >> 1) - 1) ] };
    bins McuDramVddLoLvRxCalib                                        = { [ (('h40010338 - 'h40000000) >> 1) : ((('h40010338 - 'h40000000 + 'd66) >> 1) - 1) ] };
    bins McuNvmFixSlimLdoForWkup                                      = { [ (('h40010354 - 'h40000000) >> 1) : ((('h40010354 - 'h40000000 + 'd10) >> 1) - 1) ] };
    bins McuDramVddAdbFromWkup                                        = { [ (('h40010360 - 'h40000000) >> 1) : ((('h40010360 - 'h40000000 + 'd472) >> 1) - 1) ] };
    bins McuDramVddLoLvTxCalib                                        = { [ (('h40010380 - 'h40000000) >> 1) : ((('h40010380 - 'h40000000 + 'd68) >> 1) - 1) ] };
    bins McuDramVddVregFllCalib                                       = { [ (('h400103c8 - 'h40000000) >> 1) : ((('h400103c8 - 'h40000000 + 'd56) >> 1) - 1) ] };
    bins McuDramActiveCharacterization                                = { [ (('h40010400 - 'h40000000) >> 1) : ((('h40010400 - 'h40000000 + 'd264) >> 1) - 1) ] };
    bins McuDramVddVregLoHv750Calib                                   = { [ (('h40010400 - 'h40000000) >> 1) : ((('h40010400 - 'h40000000 + 'd56) >> 1) - 1) ] };
    bins McuDramVddLcAuxCalib                                         = { [ (('h40010438 - 'h40000000) >> 1) : ((('h40010438 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins McuDramVddTempSensCalib                                      = { [ (('h40010478 - 'h40000000) >> 1) : ((('h40010478 - 'h40000000 + 'd58) >> 1) - 1) ] };
    bins vdd_adb_trim                                                 = { [ (('h400104b4 - 'h40000000) >> 1) : ((('h400104b4 - 'h40000000 + 'd12) >> 1) - 1) ] };
    bins vdd_dig_trim                                                 = { [ (('h400104c0 - 'h40000000) >> 1) : ((('h400104c0 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins vdd_sym_600_trim                                             = { [ (('h400104d0 - 'h40000000) >> 1) : ((('h400104d0 - 'h40000000 + 'd7) >> 1) - 1) ] };
    bins vdd_sym_750_trim                                             = { [ (('h400104d8 - 'h40000000) >> 1) : ((('h400104d8 - 'h40000000 + 'd8) >> 1) - 1) ] };
    bins vdd_cbias_525_trim                                           = { [ (('h400104e0 - 'h40000000) >> 1) : ((('h400104e0 - 'h40000000 + 'd7) >> 1) - 1) ] };
    bins vdd_cbias_175_trim                                           = { [ (('h400104e8 - 'h40000000) >> 1) : ((('h400104e8 - 'h40000000 + 'd32) >> 1) - 1) ] };
    bins McuDramRtcCharacterization                                   = { [ (('h40010508 - 'h40000000) >> 1) : ((('h40010508 - 'h40000000 + 'd318) >> 1) - 1) ] };
    bins vdd_lolv_trim                                                = { [ (('h40010508 - 'h40000000) >> 1) : ((('h40010508 - 'h40000000 + 'd8) >> 1) - 1) ] };
    bins vdd_vreg_fll_trim                                            = { [ (('h40010510 - 'h40000000) >> 1) : ((('h40010510 - 'h40000000 + 'd12) >> 1) - 1) ] };
    bins vdd_vreg_lohv_750_trim                                       = { [ (('h4001051c - 'h40000000) >> 1) : ((('h4001051c - 'h40000000 + 'd8) >> 1) - 1) ] };
    bins vdd_lc_aux_trim                                              = { [ (('h40010524 - 'h40000000) >> 1) : ((('h40010524 - 'h40000000 + 'd12) >> 1) - 1) ] };
    bins vdd_temp_sens_trim                                           = { [ (('h40010530 - 'h40000000) >> 1) : ((('h40010530 - 'h40000000 + 'd8) >> 1) - 1) ] };
    bins dram_vdd_adb_trim                                            = { [ (('h40010538 - 'h40000000) >> 1) : ((('h40010538 - 'h40000000 + 'd12) >> 1) - 1) ] };
    bins McuDramConfigGnvmForFllTdcCalib                              = { [ (('h40010588 - 'h40000000) >> 1) : ((('h40010588 - 'h40000000 + 'd160) >> 1) - 1) ] };
    bins McuNvmTurnOnTdcAndSetFirstTrim                               = { [ (('h40010628 - 'h40000000) >> 1) : ((('h40010628 - 'h40000000 + 'd40) >> 1) - 1) ] };
    bins rtc_clk_char_trim_dram                                       = { [ (('h40010648 - 'h40000000) >> 1) : ((('h40010648 - 'h40000000 + 'd16) >> 1) - 1) ] };
    bins vstart_trim_nvm                                              = { [ (('h40010650 - 'h40000000) >> 1) : ((('h40010650 - 'h40000000 + 'd128) >> 1) - 1) ] };